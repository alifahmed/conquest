module conquest_tb();

    // Generated top module signals
    reg  clk_i;
    reg  rst_i;
    reg  [31:0] m0_data_i = 32'b0;
    wire [31:0] m0_data_o;
    reg  [31:0] m0_addr_i = 32'b0;
    reg  [3:0] m0_sel_i = 4'b0;
    reg  m0_we_i = 1'b0;
    reg  m0_cyc_i = 1'b0;
    reg  m0_stb_i = 1'b0;
    wire m0_ack_o;
    wire m0_err_o;
    wire m0_rty_o;
    reg  [31:0] m1_data_i = 32'b0;
    wire [31:0] m1_data_o;
    reg  [31:0] m1_addr_i = 32'b0;
    reg  [3:0] m1_sel_i = 4'b0;
    reg  m1_we_i = 1'b0;
    reg  m1_cyc_i = 1'b0;
    reg  m1_stb_i = 1'b0;
    wire m1_ack_o;
    wire m1_err_o;
    wire m1_rty_o;
    reg  [31:0] m2_data_i = 32'b0;
    wire [31:0] m2_data_o;
    reg  [31:0] m2_addr_i = 32'b0;
    reg  [3:0] m2_sel_i = 4'b0;
    reg  m2_we_i = 1'b0;
    reg  m2_cyc_i = 1'b0;
    reg  m2_stb_i = 1'b0;
    wire m2_ack_o;
    wire m2_err_o;
    wire m2_rty_o;
    reg  [31:0] m3_data_i = 32'b0;
    wire [31:0] m3_data_o;
    reg  [31:0] m3_addr_i = 32'b0;
    reg  [3:0] m3_sel_i = 4'b0;
    reg  m3_we_i = 1'b0;
    reg  m3_cyc_i = 1'b0;
    reg  m3_stb_i = 1'b0;
    wire m3_ack_o;
    wire m3_err_o;
    wire m3_rty_o;
    reg  [31:0] m4_data_i = 32'b0;
    wire [31:0] m4_data_o;
    reg  [31:0] m4_addr_i = 32'b0;
    reg  [3:0] m4_sel_i = 4'b0;
    reg  m4_we_i = 1'b0;
    reg  m4_cyc_i = 1'b0;
    reg  m4_stb_i = 1'b0;
    wire m4_ack_o;
    wire m4_err_o;
    wire m4_rty_o;
    reg  [31:0] m5_data_i = 32'b0;
    wire [31:0] m5_data_o;
    reg  [31:0] m5_addr_i = 32'b0;
    reg  [3:0] m5_sel_i = 4'b0;
    reg  m5_we_i = 1'b0;
    reg  m5_cyc_i = 1'b0;
    reg  m5_stb_i = 1'b0;
    wire m5_ack_o;
    wire m5_err_o;
    wire m5_rty_o;
    reg  [31:0] m6_data_i = 32'b0;
    wire [31:0] m6_data_o;
    reg  [31:0] m6_addr_i = 32'b0;
    reg  [3:0] m6_sel_i = 4'b0;
    reg  m6_we_i = 1'b0;
    reg  m6_cyc_i = 1'b0;
    reg  m6_stb_i = 1'b0;
    wire m6_ack_o;
    wire m6_err_o;
    wire m6_rty_o;
    reg  [31:0] m7_data_i = 32'b0;
    wire [31:0] m7_data_o;
    reg  [31:0] m7_addr_i = 32'b0;
    reg  [3:0] m7_sel_i = 4'b0;
    reg  m7_we_i = 1'b0;
    reg  m7_cyc_i = 1'b0;
    reg  m7_stb_i = 1'b0;
    wire m7_ack_o;
    wire m7_err_o;
    wire m7_rty_o;
    reg  [31:0] s0_data_i = 32'b0;
    wire [31:0] s0_data_o;
    wire [31:0] s0_addr_o;
    wire [3:0] s0_sel_o;
    wire s0_we_o;
    wire s0_cyc_o;
    wire s0_stb_o;
    reg  s0_ack_i = 1'b0;
    reg  s0_err_i = 1'b0;
    reg  s0_rty_i = 1'b0;
    reg  [31:0] s1_data_i = 32'b0;
    wire [31:0] s1_data_o;
    wire [31:0] s1_addr_o;
    wire [3:0] s1_sel_o;
    wire s1_we_o;
    wire s1_cyc_o;
    wire s1_stb_o;
    reg  s1_ack_i = 1'b0;
    reg  s1_err_i = 1'b0;
    reg  s1_rty_i = 1'b0;
    reg  [31:0] s2_data_i = 32'b0;
    wire [31:0] s2_data_o;
    wire [31:0] s2_addr_o;
    wire [3:0] s2_sel_o;
    wire s2_we_o;
    wire s2_cyc_o;
    wire s2_stb_o;
    reg  s2_ack_i = 1'b0;
    reg  s2_err_i = 1'b0;
    reg  s2_rty_i = 1'b0;
    reg  [31:0] s3_data_i = 32'b0;
    wire [31:0] s3_data_o;
    wire [31:0] s3_addr_o;
    wire [3:0] s3_sel_o;
    wire s3_we_o;
    wire s3_cyc_o;
    wire s3_stb_o;
    reg  s3_ack_i = 1'b0;
    reg  s3_err_i = 1'b0;
    reg  s3_rty_i = 1'b0;
    reg  [31:0] s4_data_i = 32'b0;
    wire [31:0] s4_data_o;
    wire [31:0] s4_addr_o;
    wire [3:0] s4_sel_o;
    wire s4_we_o;
    wire s4_cyc_o;
    wire s4_stb_o;
    reg  s4_ack_i = 1'b0;
    reg  s4_err_i = 1'b0;
    reg  s4_rty_i = 1'b0;
    reg  [31:0] s5_data_i = 32'b0;
    wire [31:0] s5_data_o;
    wire [31:0] s5_addr_o;
    wire [3:0] s5_sel_o;
    wire s5_we_o;
    wire s5_cyc_o;
    wire s5_stb_o;
    reg  s5_ack_i = 1'b0;
    reg  s5_err_i = 1'b0;
    reg  s5_rty_i = 1'b0;
    reg  [31:0] s6_data_i = 32'b0;
    wire [31:0] s6_data_o;
    wire [31:0] s6_addr_o;
    wire [3:0] s6_sel_o;
    wire s6_we_o;
    wire s6_cyc_o;
    wire s6_stb_o;
    reg  s6_ack_i = 1'b0;
    reg  s6_err_i = 1'b0;
    reg  s6_rty_i = 1'b0;
    reg  [31:0] s7_data_i = 32'b0;
    wire [31:0] s7_data_o;
    wire [31:0] s7_addr_o;
    wire [3:0] s7_sel_o;
    wire s7_we_o;
    wire s7_cyc_o;
    wire s7_stb_o;
    reg  s7_ack_i = 1'b0;
    reg  s7_err_i = 1'b0;
    reg  s7_rty_i = 1'b0;
    reg  [31:0] s8_data_i = 32'b0;
    wire [31:0] s8_data_o;
    wire [31:0] s8_addr_o;
    wire [3:0] s8_sel_o;
    wire s8_we_o;
    wire s8_cyc_o;
    wire s8_stb_o;
    reg  s8_ack_i = 1'b0;
    reg  s8_err_i = 1'b0;
    reg  s8_rty_i = 1'b0;
    reg  [31:0] s9_data_i = 32'b0;
    wire [31:0] s9_data_o;
    wire [31:0] s9_addr_o;
    wire [3:0] s9_sel_o;
    wire s9_we_o;
    wire s9_cyc_o;
    wire s9_stb_o;
    reg  s9_ack_i = 1'b0;
    reg  s9_err_i = 1'b0;
    reg  s9_rty_i = 1'b0;
    reg  [31:0] s10_data_i = 32'b0;
    wire [31:0] s10_data_o;
    wire [31:0] s10_addr_o;
    wire [3:0] s10_sel_o;
    wire s10_we_o;
    wire s10_cyc_o;
    wire s10_stb_o;
    reg  s10_ack_i = 1'b0;
    reg  s10_err_i = 1'b0;
    reg  s10_rty_i = 1'b0;
    reg  [31:0] s11_data_i = 32'b0;
    wire [31:0] s11_data_o;
    wire [31:0] s11_addr_o;
    wire [3:0] s11_sel_o;
    wire s11_we_o;
    wire s11_cyc_o;
    wire s11_stb_o;
    reg  s11_ack_i = 1'b0;
    reg  s11_err_i = 1'b0;
    reg  s11_rty_i = 1'b0;
    reg  [31:0] s12_data_i = 32'b0;
    wire [31:0] s12_data_o;
    wire [31:0] s12_addr_o;
    wire [3:0] s12_sel_o;
    wire s12_we_o;
    wire s12_cyc_o;
    wire s12_stb_o;
    reg  s12_ack_i = 1'b0;
    reg  s12_err_i = 1'b0;
    reg  s12_rty_i = 1'b0;
    reg  [31:0] s13_data_i = 32'b0;
    wire [31:0] s13_data_o;
    wire [31:0] s13_addr_o;
    wire [3:0] s13_sel_o;
    wire s13_we_o;
    wire s13_cyc_o;
    wire s13_stb_o;
    reg  s13_ack_i = 1'b0;
    reg  s13_err_i = 1'b0;
    reg  s13_rty_i = 1'b0;
    reg  [31:0] s14_data_i = 32'b0;
    wire [31:0] s14_data_o;
    wire [31:0] s14_addr_o;
    wire [3:0] s14_sel_o;
    wire s14_we_o;
    wire s14_cyc_o;
    wire s14_stb_o;
    reg  s14_ack_i = 1'b0;
    reg  s14_err_i = 1'b0;
    reg  s14_rty_i = 1'b0;
    reg  [31:0] s15_data_i = 32'b0;
    wire [31:0] s15_data_o;
    wire [31:0] s15_addr_o;
    wire [3:0] s15_sel_o;
    wire s15_we_o;
    wire s15_cyc_o;
    wire s15_stb_o;
    reg  s15_ack_i = 1'b0;
    reg  s15_err_i = 1'b0;
    reg  s15_rty_i = 1'b0;
    reg  __obs;

    // Generated top module instance
    wb_conmax_top _conc_top_inst(
            .clk_i     ( clk_i ),
            .rst_i     ( rst_i ),
            .m0_data_i ( m0_data_i ),
            .m0_data_o ( m0_data_o ),
            .m0_addr_i ( m0_addr_i ),
            .m0_sel_i  ( m0_sel_i ),
            .m0_we_i   ( m0_we_i ),
            .m0_cyc_i  ( m0_cyc_i ),
            .m0_stb_i  ( m0_stb_i ),
            .m0_ack_o  ( m0_ack_o ),
            .m0_err_o  ( m0_err_o ),
            .m0_rty_o  ( m0_rty_o ),
            .m1_data_i ( m1_data_i ),
            .m1_data_o ( m1_data_o ),
            .m1_addr_i ( m1_addr_i ),
            .m1_sel_i  ( m1_sel_i ),
            .m1_we_i   ( m1_we_i ),
            .m1_cyc_i  ( m1_cyc_i ),
            .m1_stb_i  ( m1_stb_i ),
            .m1_ack_o  ( m1_ack_o ),
            .m1_err_o  ( m1_err_o ),
            .m1_rty_o  ( m1_rty_o ),
            .m2_data_i ( m2_data_i ),
            .m2_data_o ( m2_data_o ),
            .m2_addr_i ( m2_addr_i ),
            .m2_sel_i  ( m2_sel_i ),
            .m2_we_i   ( m2_we_i ),
            .m2_cyc_i  ( m2_cyc_i ),
            .m2_stb_i  ( m2_stb_i ),
            .m2_ack_o  ( m2_ack_o ),
            .m2_err_o  ( m2_err_o ),
            .m2_rty_o  ( m2_rty_o ),
            .m3_data_i ( m3_data_i ),
            .m3_data_o ( m3_data_o ),
            .m3_addr_i ( m3_addr_i ),
            .m3_sel_i  ( m3_sel_i ),
            .m3_we_i   ( m3_we_i ),
            .m3_cyc_i  ( m3_cyc_i ),
            .m3_stb_i  ( m3_stb_i ),
            .m3_ack_o  ( m3_ack_o ),
            .m3_err_o  ( m3_err_o ),
            .m3_rty_o  ( m3_rty_o ),
            .m4_data_i ( m4_data_i ),
            .m4_data_o ( m4_data_o ),
            .m4_addr_i ( m4_addr_i ),
            .m4_sel_i  ( m4_sel_i ),
            .m4_we_i   ( m4_we_i ),
            .m4_cyc_i  ( m4_cyc_i ),
            .m4_stb_i  ( m4_stb_i ),
            .m4_ack_o  ( m4_ack_o ),
            .m4_err_o  ( m4_err_o ),
            .m4_rty_o  ( m4_rty_o ),
            .m5_data_i ( m5_data_i ),
            .m5_data_o ( m5_data_o ),
            .m5_addr_i ( m5_addr_i ),
            .m5_sel_i  ( m5_sel_i ),
            .m5_we_i   ( m5_we_i ),
            .m5_cyc_i  ( m5_cyc_i ),
            .m5_stb_i  ( m5_stb_i ),
            .m5_ack_o  ( m5_ack_o ),
            .m5_err_o  ( m5_err_o ),
            .m5_rty_o  ( m5_rty_o ),
            .m6_data_i ( m6_data_i ),
            .m6_data_o ( m6_data_o ),
            .m6_addr_i ( m6_addr_i ),
            .m6_sel_i  ( m6_sel_i ),
            .m6_we_i   ( m6_we_i ),
            .m6_cyc_i  ( m6_cyc_i ),
            .m6_stb_i  ( m6_stb_i ),
            .m6_ack_o  ( m6_ack_o ),
            .m6_err_o  ( m6_err_o ),
            .m6_rty_o  ( m6_rty_o ),
            .m7_data_i ( m7_data_i ),
            .m7_data_o ( m7_data_o ),
            .m7_addr_i ( m7_addr_i ),
            .m7_sel_i  ( m7_sel_i ),
            .m7_we_i   ( m7_we_i ),
            .m7_cyc_i  ( m7_cyc_i ),
            .m7_stb_i  ( m7_stb_i ),
            .m7_ack_o  ( m7_ack_o ),
            .m7_err_o  ( m7_err_o ),
            .m7_rty_o  ( m7_rty_o ),
            .s0_data_i ( s0_data_i ),
            .s0_data_o ( s0_data_o ),
            .s0_addr_o ( s0_addr_o ),
            .s0_sel_o  ( s0_sel_o ),
            .s0_we_o   ( s0_we_o ),
            .s0_cyc_o  ( s0_cyc_o ),
            .s0_stb_o  ( s0_stb_o ),
            .s0_ack_i  ( s0_ack_i ),
            .s0_err_i  ( s0_err_i ),
            .s0_rty_i  ( s0_rty_i ),
            .s1_data_i ( s1_data_i ),
            .s1_data_o ( s1_data_o ),
            .s1_addr_o ( s1_addr_o ),
            .s1_sel_o  ( s1_sel_o ),
            .s1_we_o   ( s1_we_o ),
            .s1_cyc_o  ( s1_cyc_o ),
            .s1_stb_o  ( s1_stb_o ),
            .s1_ack_i  ( s1_ack_i ),
            .s1_err_i  ( s1_err_i ),
            .s1_rty_i  ( s1_rty_i ),
            .s2_data_i ( s2_data_i ),
            .s2_data_o ( s2_data_o ),
            .s2_addr_o ( s2_addr_o ),
            .s2_sel_o  ( s2_sel_o ),
            .s2_we_o   ( s2_we_o ),
            .s2_cyc_o  ( s2_cyc_o ),
            .s2_stb_o  ( s2_stb_o ),
            .s2_ack_i  ( s2_ack_i ),
            .s2_err_i  ( s2_err_i ),
            .s2_rty_i  ( s2_rty_i ),
            .s3_data_i ( s3_data_i ),
            .s3_data_o ( s3_data_o ),
            .s3_addr_o ( s3_addr_o ),
            .s3_sel_o  ( s3_sel_o ),
            .s3_we_o   ( s3_we_o ),
            .s3_cyc_o  ( s3_cyc_o ),
            .s3_stb_o  ( s3_stb_o ),
            .s3_ack_i  ( s3_ack_i ),
            .s3_err_i  ( s3_err_i ),
            .s3_rty_i  ( s3_rty_i ),
            .s4_data_i ( s4_data_i ),
            .s4_data_o ( s4_data_o ),
            .s4_addr_o ( s4_addr_o ),
            .s4_sel_o  ( s4_sel_o ),
            .s4_we_o   ( s4_we_o ),
            .s4_cyc_o  ( s4_cyc_o ),
            .s4_stb_o  ( s4_stb_o ),
            .s4_ack_i  ( s4_ack_i ),
            .s4_err_i  ( s4_err_i ),
            .s4_rty_i  ( s4_rty_i ),
            .s5_data_i ( s5_data_i ),
            .s5_data_o ( s5_data_o ),
            .s5_addr_o ( s5_addr_o ),
            .s5_sel_o  ( s5_sel_o ),
            .s5_we_o   ( s5_we_o ),
            .s5_cyc_o  ( s5_cyc_o ),
            .s5_stb_o  ( s5_stb_o ),
            .s5_ack_i  ( s5_ack_i ),
            .s5_err_i  ( s5_err_i ),
            .s5_rty_i  ( s5_rty_i ),
            .s6_data_i ( s6_data_i ),
            .s6_data_o ( s6_data_o ),
            .s6_addr_o ( s6_addr_o ),
            .s6_sel_o  ( s6_sel_o ),
            .s6_we_o   ( s6_we_o ),
            .s6_cyc_o  ( s6_cyc_o ),
            .s6_stb_o  ( s6_stb_o ),
            .s6_ack_i  ( s6_ack_i ),
            .s6_err_i  ( s6_err_i ),
            .s6_rty_i  ( s6_rty_i ),
            .s7_data_i ( s7_data_i ),
            .s7_data_o ( s7_data_o ),
            .s7_addr_o ( s7_addr_o ),
            .s7_sel_o  ( s7_sel_o ),
            .s7_we_o   ( s7_we_o ),
            .s7_cyc_o  ( s7_cyc_o ),
            .s7_stb_o  ( s7_stb_o ),
            .s7_ack_i  ( s7_ack_i ),
            .s7_err_i  ( s7_err_i ),
            .s7_rty_i  ( s7_rty_i ),
            .s8_data_i ( s8_data_i ),
            .s8_data_o ( s8_data_o ),
            .s8_addr_o ( s8_addr_o ),
            .s8_sel_o  ( s8_sel_o ),
            .s8_we_o   ( s8_we_o ),
            .s8_cyc_o  ( s8_cyc_o ),
            .s8_stb_o  ( s8_stb_o ),
            .s8_ack_i  ( s8_ack_i ),
            .s8_err_i  ( s8_err_i ),
            .s8_rty_i  ( s8_rty_i ),
            .s9_data_i ( s9_data_i ),
            .s9_data_o ( s9_data_o ),
            .s9_addr_o ( s9_addr_o ),
            .s9_sel_o  ( s9_sel_o ),
            .s9_we_o   ( s9_we_o ),
            .s9_cyc_o  ( s9_cyc_o ),
            .s9_stb_o  ( s9_stb_o ),
            .s9_ack_i  ( s9_ack_i ),
            .s9_err_i  ( s9_err_i ),
            .s9_rty_i  ( s9_rty_i ),
            .s10_data_i( s10_data_i ),
            .s10_data_o( s10_data_o ),
            .s10_addr_o( s10_addr_o ),
            .s10_sel_o ( s10_sel_o ),
            .s10_we_o  ( s10_we_o ),
            .s10_cyc_o ( s10_cyc_o ),
            .s10_stb_o ( s10_stb_o ),
            .s10_ack_i ( s10_ack_i ),
            .s10_err_i ( s10_err_i ),
            .s10_rty_i ( s10_rty_i ),
            .s11_data_i( s11_data_i ),
            .s11_data_o( s11_data_o ),
            .s11_addr_o( s11_addr_o ),
            .s11_sel_o ( s11_sel_o ),
            .s11_we_o  ( s11_we_o ),
            .s11_cyc_o ( s11_cyc_o ),
            .s11_stb_o ( s11_stb_o ),
            .s11_ack_i ( s11_ack_i ),
            .s11_err_i ( s11_err_i ),
            .s11_rty_i ( s11_rty_i ),
            .s12_data_i( s12_data_i ),
            .s12_data_o( s12_data_o ),
            .s12_addr_o( s12_addr_o ),
            .s12_sel_o ( s12_sel_o ),
            .s12_we_o  ( s12_we_o ),
            .s12_cyc_o ( s12_cyc_o ),
            .s12_stb_o ( s12_stb_o ),
            .s12_ack_i ( s12_ack_i ),
            .s12_err_i ( s12_err_i ),
            .s12_rty_i ( s12_rty_i ),
            .s13_data_i( s13_data_i ),
            .s13_data_o( s13_data_o ),
            .s13_addr_o( s13_addr_o ),
            .s13_sel_o ( s13_sel_o ),
            .s13_we_o  ( s13_we_o ),
            .s13_cyc_o ( s13_cyc_o ),
            .s13_stb_o ( s13_stb_o ),
            .s13_ack_i ( s13_ack_i ),
            .s13_err_i ( s13_err_i ),
            .s13_rty_i ( s13_rty_i ),
            .s14_data_i( s14_data_i ),
            .s14_data_o( s14_data_o ),
            .s14_addr_o( s14_addr_o ),
            .s14_sel_o ( s14_sel_o ),
            .s14_we_o  ( s14_we_o ),
            .s14_cyc_o ( s14_cyc_o ),
            .s14_stb_o ( s14_stb_o ),
            .s14_ack_i ( s14_ack_i ),
            .s14_err_i ( s14_err_i ),
            .s14_rty_i ( s14_rty_i ),
            .s15_data_i( s15_data_i ),
            .s15_data_o( s15_data_o ),
            .s15_addr_o( s15_addr_o ),
            .s15_sel_o ( s15_sel_o ),
            .s15_we_o  ( s15_we_o ),
            .s15_cyc_o ( s15_cyc_o ),
            .s15_stb_o ( s15_stb_o ),
            .s15_ack_i ( s15_ack_i ),
            .s15_err_i ( s15_err_i ),
            .s15_rty_i ( s15_rty_i ),
            .__obs     ( __obs ));

    // Generated internal use signals
    reg  [31:0] _conc_pc;
    reg  [1128:0] _conc_opcode;
    reg  [1128:0] _conc_ram[0:10];


    // Generated clock pulse
    always begin
        #5 clk_i = ~clk_i;
    end

    // Generated program counter
    always @(posedge clk_i) begin
        _conc_pc = _conc_pc + 32'b1;
        _conc_opcode = _conc_ram[_conc_pc];
        __obs <= #1 _conc_opcode[1128];
        m0_addr_i <= #1 _conc_opcode[63:32];
        m0_cyc_i <= #1 _conc_opcode[69];
        m0_data_i <= #1 _conc_opcode[31:0];
        m0_sel_i <= #1 _conc_opcode[67:64];
        m0_stb_i <= #1 _conc_opcode[70];
        m0_we_i <= #1 _conc_opcode[68];
        m1_addr_i <= #1 _conc_opcode[134:103];
        m1_cyc_i <= #1 _conc_opcode[140];
        m1_data_i <= #1 _conc_opcode[102:71];
        m1_sel_i <= #1 _conc_opcode[138:135];
        m1_stb_i <= #1 _conc_opcode[141];
        m1_we_i <= #1 _conc_opcode[139];
        m2_addr_i <= #1 _conc_opcode[205:174];
        m2_cyc_i <= #1 _conc_opcode[211];
        m2_data_i <= #1 _conc_opcode[173:142];
        m2_sel_i <= #1 _conc_opcode[209:206];
        m2_stb_i <= #1 _conc_opcode[212];
        m2_we_i <= #1 _conc_opcode[210];
        m3_addr_i <= #1 _conc_opcode[276:245];
        m3_cyc_i <= #1 _conc_opcode[282];
        m3_data_i <= #1 _conc_opcode[244:213];
        m3_sel_i <= #1 _conc_opcode[280:277];
        m3_stb_i <= #1 _conc_opcode[283];
        m3_we_i <= #1 _conc_opcode[281];
        m4_addr_i <= #1 _conc_opcode[347:316];
        m4_cyc_i <= #1 _conc_opcode[353];
        m4_data_i <= #1 _conc_opcode[315:284];
        m4_sel_i <= #1 _conc_opcode[351:348];
        m4_stb_i <= #1 _conc_opcode[354];
        m4_we_i <= #1 _conc_opcode[352];
        m5_addr_i <= #1 _conc_opcode[418:387];
        m5_cyc_i <= #1 _conc_opcode[424];
        m5_data_i <= #1 _conc_opcode[386:355];
        m5_sel_i <= #1 _conc_opcode[422:419];
        m5_stb_i <= #1 _conc_opcode[425];
        m5_we_i <= #1 _conc_opcode[423];
        m6_addr_i <= #1 _conc_opcode[489:458];
        m6_cyc_i <= #1 _conc_opcode[495];
        m6_data_i <= #1 _conc_opcode[457:426];
        m6_sel_i <= #1 _conc_opcode[493:490];
        m6_stb_i <= #1 _conc_opcode[496];
        m6_we_i <= #1 _conc_opcode[494];
        m7_addr_i <= #1 _conc_opcode[560:529];
        m7_cyc_i <= #1 _conc_opcode[566];
        m7_data_i <= #1 _conc_opcode[528:497];
        m7_sel_i <= #1 _conc_opcode[564:561];
        m7_stb_i <= #1 _conc_opcode[567];
        m7_we_i <= #1 _conc_opcode[565];
        s0_ack_i <= #1 _conc_opcode[600];
        s0_data_i <= #1 _conc_opcode[599:568];
        s0_err_i <= #1 _conc_opcode[601];
        s0_rty_i <= #1 _conc_opcode[602];
        s10_ack_i <= #1 _conc_opcode[950];
        s10_data_i <= #1 _conc_opcode[949:918];
        s10_err_i <= #1 _conc_opcode[951];
        s10_rty_i <= #1 _conc_opcode[952];
        s11_ack_i <= #1 _conc_opcode[985];
        s11_data_i <= #1 _conc_opcode[984:953];
        s11_err_i <= #1 _conc_opcode[986];
        s11_rty_i <= #1 _conc_opcode[987];
        s12_ack_i <= #1 _conc_opcode[1020];
        s12_data_i <= #1 _conc_opcode[1019:988];
        s12_err_i <= #1 _conc_opcode[1021];
        s12_rty_i <= #1 _conc_opcode[1022];
        s13_ack_i <= #1 _conc_opcode[1055];
        s13_data_i <= #1 _conc_opcode[1054:1023];
        s13_err_i <= #1 _conc_opcode[1056];
        s13_rty_i <= #1 _conc_opcode[1057];
        s14_ack_i <= #1 _conc_opcode[1090];
        s14_data_i <= #1 _conc_opcode[1089:1058];
        s14_err_i <= #1 _conc_opcode[1091];
        s14_rty_i <= #1 _conc_opcode[1092];
        s15_ack_i <= #1 _conc_opcode[1125];
        s15_data_i <= #1 _conc_opcode[1124:1093];
        s15_err_i <= #1 _conc_opcode[1126];
        s15_rty_i <= #1 _conc_opcode[1127];
        s1_ack_i <= #1 _conc_opcode[635];
        s1_data_i <= #1 _conc_opcode[634:603];
        s1_err_i <= #1 _conc_opcode[636];
        s1_rty_i <= #1 _conc_opcode[637];
        s2_ack_i <= #1 _conc_opcode[670];
        s2_data_i <= #1 _conc_opcode[669:638];
        s2_err_i <= #1 _conc_opcode[671];
        s2_rty_i <= #1 _conc_opcode[672];
        s3_ack_i <= #1 _conc_opcode[705];
        s3_data_i <= #1 _conc_opcode[704:673];
        s3_err_i <= #1 _conc_opcode[706];
        s3_rty_i <= #1 _conc_opcode[707];
        s4_ack_i <= #1 _conc_opcode[740];
        s4_data_i <= #1 _conc_opcode[739:708];
        s4_err_i <= #1 _conc_opcode[741];
        s4_rty_i <= #1 _conc_opcode[742];
        s5_ack_i <= #1 _conc_opcode[775];
        s5_data_i <= #1 _conc_opcode[774:743];
        s5_err_i <= #1 _conc_opcode[776];
        s5_rty_i <= #1 _conc_opcode[777];
        s6_ack_i <= #1 _conc_opcode[810];
        s6_data_i <= #1 _conc_opcode[809:778];
        s6_err_i <= #1 _conc_opcode[811];
        s6_rty_i <= #1 _conc_opcode[812];
        s7_ack_i <= #1 _conc_opcode[845];
        s7_data_i <= #1 _conc_opcode[844:813];
        s7_err_i <= #1 _conc_opcode[846];
        s7_rty_i <= #1 _conc_opcode[847];
        s8_ack_i <= #1 _conc_opcode[880];
        s8_data_i <= #1 _conc_opcode[879:848];
        s8_err_i <= #1 _conc_opcode[881];
        s8_rty_i <= #1 _conc_opcode[882];
        s9_ack_i <= #1 _conc_opcode[915];
        s9_data_i <= #1 _conc_opcode[914:883];
        s9_err_i <= #1 _conc_opcode[916];
        s9_rty_i <= #1 _conc_opcode[917];
        $strobe(";_C %d", _conc_pc);
    end

    // Generated initial block
    initial begin
        clk_i = 1'b0;
        rst_i = 1'b0;
        _conc_pc = 32'b0;
        $readmemb("data.mem", _conc_ram);
        #2 clk_i = 1'b1;
        rst_i = 1'b1;
        #5 rst_i = 1'b0;
        #100 $finish;
    end

endmodule
