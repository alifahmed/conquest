// Following code segment is generated from ./src/b14.v:16
module b14(clock, reset, datai, addr, datao, rd, wr, __obs);
    input clock;
    input reset;
    input [30:0] datai;
    output [19:0] addr;
    output [30:0] datao;
    output rd;
    output wr;
    input __obs;

    reg B = 1'b0;
    reg [30:0] IR = 31'b0;
    reg [19:0] addr = 20'b0;
    reg cf = 1'b0;
    reg [1:0] d = 2'b0;
    reg [30:0] datao = 31'b0;
    reg [2:0] df = 3'b0;
    reg [3:0] ff = 4'b0;
    reg [30:0] m = 31'b0;
    reg [1:0] mf = 2'b0;
    reg rd = 1'b0;
    reg [30:0] reg0 = 31'b0;
    reg [30:0] reg1 = 31'b0;
    reg [30:0] reg2 = 31'b0;
    reg [30:0] reg3 = 31'b0;
    reg [30:0] rx = 31'b0;
    reg [1:0] s = 2'b0;
    reg state = 1'b0;
    reg [30:0] t = 31'b0;
    reg [19:0] tail = 20'b0;
    reg wr = 1'b0;

    always @(*) begin
        mf = IR[28:27]; $display(";A 0");		//(assert (= @mf    (bv-extract 28 27 #IR ))) ;0 BL
    end

    always @(*) begin
        df = IR[26:24]; $display(";A 1");		//(assert (= @df    (bv-extract 26 24 #IR ))) ;1 BL
    end

    always @(*) begin
        ff = IR[22:19]; $display(";A 2");		//(assert (= @ff    (bv-extract 22 19 #IR ))) ;2 BL
    end

    always @(*) begin
        cf = IR[23]; $display(";A 3");		//(assert (= @cf    (bv-extract 23 23 #IR ))) ;3 BL
    end

    always @(*) begin
        tail = IR[19:0]; $display(";A 4");		//(assert (= @tail    (bv-extract 19 0 #IR ))) ;4 BL
    end

    always @(*) begin
        s = IR[30:29]; $display(";A 5");		//(assert (= @s    (bv-extract 30 29 #IR ))) ;5 BL
    end

    // Following code segment is generated from ./src/b14.v:72
    always @(posedge clock) begin
        if ((reset == 1'b1)) begin
            IR <= #1 31'b0000000000000000000000000000000; $display(";A 8");		//(assert (= @IR    0b0000000000000000000000000000000)) ;8 NB
            d <= #1 2'b00; $display(";A 9");		//(assert (= @d    0b00)) ;9 NB
            rx <= #1 31'b0000000000000000000000000000000; $display(";A 10");		//(assert (= @rx    0b0000000000000000000000000000000)) ;10 NB
            m <= #1 31'b0000000000000000000000000000000; $display(";A 11");		//(assert (= @m    0b0000000000000000000000000000000)) ;11 NB
            B <= #1 1'b0; $display(";A 12");		//(assert (= @B    0b0)) ;12 NB
            reg0 <= #1 31'b0000000000000000000000000000000; $display(";A 13");		//(assert (= @reg0    0b0000000000000000000000000000000)) ;13 NB
            reg1 <= #1 31'b0000000000000000000000000000000; $display(";A 14");		//(assert (= @reg1    0b0000000000000000000000000000000)) ;14 NB
            reg2 <= #1 31'b0000000000000000000000000000000; $display(";A 15");		//(assert (= @reg2    0b0000000000000000000000000000000)) ;15 NB
            reg3 <= #1 31'b0000000000000000000000000000000; $display(";A 16");		//(assert (= @reg3    0b0000000000000000000000000000000)) ;16 NB
            addr <= #1 20'b00000000000000000000; $display(";A 17");		//(assert (= @addr    0b00000000000000000000)) ;17 NB
            rd <= #1 1'b0; $display(";A 18");		//(assert (= @rd    0b0)) ;18 NB
            wr <= #1 1'b0; $display(";A 19");		//(assert (= @wr    0b0)) ;19 NB
            datao <= #1 31'b0000000000000000000000000000000; $display(";A 20");		//(assert (= @datao    0b0000000000000000000000000000000)) ;20 NB
            state <= #1 1'b0; $display(";A 21");		//(assert (= @state    0b0)) ;21 NB
        end
        else begin
            case (state)
                1'b0 :
                    begin
                        $display(";A 22");		//(assert (= #state    0b0)) ;22 CS
                        addr <= #1 reg3[19:0]; $display(";A 23");		//(assert (= @addr    (bv-extract 19 0 #reg3 ))) ;23 NB
                        rd <= #1 1'b1; $display(";A 24");		//(assert (= @rd    0b1)) ;24 NB
                        IR <= #1 datai; $display(";A 25");		//(assert (= @IR    #datai )) ;25 NB
                        state <= #1 1'b1; $display(";A 26");		//(assert (= @state    0b1)) ;26 NB
                        case (datai[30:29])
                            2'b00 :
                                begin
                                    $display(";A 27");		//(assert (= (bv-extract 30 29 #datai )   0b00)) ;27 CS
                                    rx <= #1 reg0; $display(";A 28");		//(assert (= @rx    #reg0 )) ;28 NB
                                end
                            2'b01 :
                                begin
                                    $display(";A 29");		//(assert (= (bv-extract 30 29 #datai )   0b01)) ;29 CS
                                    rx <= #1 reg1; $display(";A 30");		//(assert (= @rx    #reg1 )) ;30 NB
                                end
                            2'b10 :
                                begin
                                    $display(";A 31");		//(assert (= (bv-extract 30 29 #datai )   0b10)) ;31 CS
                                    rx <= #1 reg2; $display(";A 32");		//(assert (= @rx    #reg2 )) ;32 NB
                                end
                            2'b11 :
                                begin
                                    $display(";A 33");		//(assert (= (bv-extract 30 29 #datai )   0b11)) ;33 CS
                                    rx <= #1 reg3; $display(";A 34");		//(assert (= @rx    #reg3 )) ;34 NB
                                end
                        endcase
                    end
                1'b1 :
                    begin
                        $display(";A 35");		//(assert (= #state    0b1)) ;35 CS
                        case (cf)
                            1'b1 :
                                begin
                                    $display(";A 36");		//(assert (= #cf    0b1)) ;36 CS
                                    case (mf)
                                        2'b00 :
                                            begin
                                                $display(";A 37");		//(assert (= #mf    0b00)) ;37 CS
                                                m = {11'b00000000000, tail}; $display(";A 38");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;38 BL
                                            end
                                        2'b01 :
                                            begin
                                                $display(";A 39");		//(assert (= #mf    0b01)) ;39 CS
                                                m = datai; $display(";A 40");		//(assert (= @m    #datai )) ;40 BL
                                                addr <= #1 tail; $display(";A 41");		//(assert (= @addr    #tail )) ;41 NB
                                                rd <= #1 1'b1; $display(";A 42");		//(assert (= @rd    0b1)) ;42 NB
                                            end
                                        2'b10 :
                                            begin
                                                $display(";A 43");		//(assert (= #mf    0b10)) ;43 CS
                                                addr <= #1 (tail + reg1[19:0]); $display(";A 44");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;44 NB
                                                rd <= #1 1'b1; $display(";A 45");		//(assert (= @rd    0b1)) ;45 NB
                                                m = datai; $display(";A 46");		//(assert (= @m    #datai )) ;46 BL
                                            end
                                        2'b11 :
                                            begin
                                                $display(";A 47");		//(assert (= #mf    0b11)) ;47 CS
                                                addr <= #1 (tail + reg2[19:0]); $display(";A 48");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;48 NB
                                                rd <= #1 1'b1; $display(";A 49");		//(assert (= @rd    0b1)) ;49 NB
                                                m = datai; $display(";A 50");		//(assert (= @m    #datai )) ;50 BL
                                            end
                                    endcase
                                    case (ff)
                                        4'b0000 :
                                            begin
                                                $display(";A 51");		//(assert (= #ff    0b0000)) ;51 CS
                                                if ((rx < m)) begin
                                                    $display(";A 52");		//(assert (= (bool-to-bv (bv-lt #rx  #m ))   0b1)) ;52 BR
                                                    B <= #1 1'b1; $display(";A 54");		//(assert (= @B    0b1)) ;54 NB
                                                end
                                                else begin
                                                    $display(";A 53");		//(assert (= (bool-to-bv (bv-lt #rx  #m ))   0b0)) ;53 BR
                                                    B <= #1 1'b0; $display(";A 55");		//(assert (= @B    0b0)) ;55 NB
                                                end
                                            end
                                        4'b0001 :
                                            begin
                                                $display(";A 56");		//(assert (= #ff    0b0001)) ;56 CS
                                                if ((rx >= m)) begin
                                                    $display(";A 57");		//(assert (= (bool-to-bv (bv-ge #rx  #m ))   0b1)) ;57 BR
                                                    B <= #1 1'b1; $display(";A 59");		//(assert (= @B    0b1)) ;59 NB
                                                end
                                                else begin
                                                    $display(";A 58");		//(assert (= (bool-to-bv (bv-ge #rx  #m ))   0b0)) ;58 BR
                                                    B <= #1 1'b0; $display(";A 60");		//(assert (= @B    0b0)) ;60 NB
                                                end
                                            end
                                        4'b0010 :
                                            begin
                                                $display(";A 61");		//(assert (= #ff    0b0010)) ;61 CS
                                                if ((rx == m)) begin
                                                    $display(";A 62");		//(assert (= (bv-comp #rx  #m )   0b1)) ;62 BR
                                                    B <= #1 1'b1; $display(";A 64");		//(assert (= @B    0b1)) ;64 NB
                                                end
                                                else begin
                                                    $display(";A 63");		//(assert (= (bv-comp #rx  #m )   0b0)) ;63 BR
                                                    B <= #1 1'b0; $display(";A 65");		//(assert (= @B    0b0)) ;65 NB
                                                end
                                            end
                                        4'b0011 :
                                            begin
                                                $display(";A 66");		//(assert (= #ff    0b0011)) ;66 CS
                                                if ((rx != m)) begin
                                                    $display(";A 67");		//(assert (= (bv-not (bv-comp #rx  #m ))   0b1)) ;67 BR
                                                    B <= #1 1'b1; $display(";A 69");		//(assert (= @B    0b1)) ;69 NB
                                                end
                                                else begin
                                                    $display(";A 68");		//(assert (= (bv-not (bv-comp #rx  #m ))   0b0)) ;68 BR
                                                    B <= #1 1'b0; $display(";A 70");		//(assert (= @B    0b0)) ;70 NB
                                                end
                                            end
                                        4'b0100 :
                                            begin
                                                $display(";A 71");		//(assert (= #ff    0b0100)) ;71 CS
                                                if ((rx <= m)) begin
                                                    $display(";A 72");		//(assert (= (bool-to-bv (bv-le #rx  #m ))   0b1)) ;72 BR
                                                    B <= #1 1'b1; $display(";A 74");		//(assert (= @B    0b1)) ;74 NB
                                                end
                                                else begin
                                                    $display(";A 73");		//(assert (= (bool-to-bv (bv-le #rx  #m ))   0b0)) ;73 BR
                                                    B <= #1 1'b0; $display(";A 75");		//(assert (= @B    0b0)) ;75 NB
                                                end
                                            end
                                        4'b0101 :
                                            begin
                                                $display(";A 76");		//(assert (= #ff    0b0101)) ;76 CS
                                                if ((rx > m)) begin
                                                    $display(";A 77");		//(assert (= (bool-to-bv (bv-gt #rx  #m ))   0b1)) ;77 BR
                                                    B <= #1 1'b1; $display(";A 79");		//(assert (= @B    0b1)) ;79 NB
                                                end
                                                else begin
                                                    $display(";A 78");		//(assert (= (bool-to-bv (bv-gt #rx  #m ))   0b0)) ;78 BR
                                                    B <= #1 1'b0; $display(";A 80");		//(assert (= @B    0b0)) ;80 NB
                                                end
                                            end
                                        4'b0110 :
                                            begin
                                                $display(";A 81");		//(assert (= #ff    0b0110)) ;81 CS
                                                if ((rx > 31'b0111111111111111111111111111111)) begin
                                                    $display(";A 82");		//(assert (= (bool-to-bv (bv-gt #rx  0b0111111111111111111111111111111))   0b1)) ;82 BR
                                                    rx = rx; $display(";A 84");		//(assert (= @rx    #rx )) ;84 BL
                                                end
                                                else begin
                                                    $display(";A 83");		//(assert (= (bool-to-bv (bv-gt #rx  0b0111111111111111111111111111111))   0b0)) ;83 BR
                                                end
                                                if ((rx < m)) begin
                                                    $display(";A 85");		//(assert (= (bool-to-bv (bv-lt #rx  #m ))   0b1)) ;85 BR
                                                    B <= #1 1'b1; $display(";A 87");		//(assert (= @B    0b1)) ;87 NB
                                                end
                                                else begin
                                                    $display(";A 86");		//(assert (= (bool-to-bv (bv-lt #rx  #m ))   0b0)) ;86 BR
                                                    B <= #1 1'b0; $display(";A 88");		//(assert (= @B    0b0)) ;88 NB
                                                end
                                            end
                                        4'b0111 :
                                            begin
                                                $display(";A 89");		//(assert (= #ff    0b0111)) ;89 CS
                                                if ((rx > 31'b0111111111111111111111111111111)) begin
                                                    $display(";A 90");		//(assert (= (bool-to-bv (bv-gt #rx  0b0111111111111111111111111111111))   0b1)) ;90 BR
                                                    rx = rx; $display(";A 92");		//(assert (= @rx    #rx )) ;92 BL
                                                end
                                                else begin
                                                    $display(";A 91");		//(assert (= (bool-to-bv (bv-gt #rx  0b0111111111111111111111111111111))   0b0)) ;91 BR
                                                end
                                                if ((rx >= m)) begin
                                                    $display(";A 93");		//(assert (= (bool-to-bv (bv-ge #rx  #m ))   0b1)) ;93 BR
                                                    B <= #1 1'b1; $display(";A 95");		//(assert (= @B    0b1)) ;95 NB
                                                end
                                                else begin
                                                    $display(";A 94");		//(assert (= (bool-to-bv (bv-ge #rx  #m ))   0b0)) ;94 BR
                                                    B <= #1 1'b0; $display(";A 96");		//(assert (= @B    0b0)) ;96 NB
                                                end
                                            end
                                        4'b1000 :
                                            begin
                                                $display(";A 97");		//(assert (= #ff    0b1000)) ;97 CS
                                                if (((rx < m) || (B == 1'b1))) begin
                                                    $display(";A 98");		//(assert (= (bv-or (bool-to-bv (bv-lt #rx  #m )) (bv-comp #B  0b1))   0b1)) ;98 BR
                                                    B <= #1 1'b1; $display(";A 100");		//(assert (= @B    0b1)) ;100 NB
                                                end
                                                else begin
                                                    $display(";A 99");		//(assert (= (bv-or (bool-to-bv (bv-lt #rx  #m )) (bv-comp #B  0b1))   0b0)) ;99 BR
                                                    B <= #1 1'b0; $display(";A 101");		//(assert (= @B    0b0)) ;101 NB
                                                end
                                            end
                                        4'b1001 :
                                            begin
                                                $display(";A 102");		//(assert (= #ff    0b1001)) ;102 CS
                                                if (((!(rx < m)) || (B == 1'b1))) begin
                                                    $display(";A 103");		//(assert (= (bv-or (bv-not (bv-redor (bool-to-bv (bv-lt #rx  #m )))) (bv-comp #B  0b1))   0b1)) ;103 BR
                                                    B <= #1 1'b1; $display(";A 105");		//(assert (= @B    0b1)) ;105 NB
                                                end
                                                else begin
                                                    $display(";A 104");		//(assert (= (bv-or (bv-not (bv-redor (bool-to-bv (bv-lt #rx  #m )))) (bv-comp #B  0b1))   0b0)) ;104 BR
                                                    B <= #1 1'b0; $display(";A 106");		//(assert (= @B    0b0)) ;106 NB
                                                end
                                            end
                                        4'b1010 :
                                            begin
                                                $display(";A 107");		//(assert (= #ff    0b1010)) ;107 CS
                                                if (((rx == m) || (B == 1'b1))) begin
                                                    $display(";A 108");		//(assert (= (bv-or (bv-comp #rx  #m ) (bv-comp #B  0b1))   0b1)) ;108 BR
                                                    B <= #1 1'b1; $display(";A 110");		//(assert (= @B    0b1)) ;110 NB
                                                end
                                                else begin
                                                    $display(";A 109");		//(assert (= (bv-or (bv-comp #rx  #m ) (bv-comp #B  0b1))   0b0)) ;109 BR
                                                    B <= #1 1'b0; $display(";A 111");		//(assert (= @B    0b0)) ;111 NB
                                                end
                                            end
                                        4'b1011 :
                                            begin
                                                $display(";A 112");		//(assert (= #ff    0b1011)) ;112 CS
                                                if (((!(rx == m)) || (B == 1'b1))) begin
                                                    $display(";A 113");		//(assert (= (bv-or (bv-not (bv-redor (bv-comp #rx  #m ))) (bv-comp #B  0b1))   0b1)) ;113 BR
                                                    B <= #1 1'b1; $display(";A 115");		//(assert (= @B    0b1)) ;115 NB
                                                end
                                                else begin
                                                    $display(";A 114");		//(assert (= (bv-or (bv-not (bv-redor (bv-comp #rx  #m ))) (bv-comp #B  0b1))   0b0)) ;114 BR
                                                    B <= #1 1'b0; $display(";A 116");		//(assert (= @B    0b0)) ;116 NB
                                                end
                                            end
                                        4'b1100 :
                                            begin
                                                $display(";A 117");		//(assert (= #ff    0b1100)) ;117 CS
                                                if (((!(rx > m)) || (B == 1'b1))) begin
                                                    $display(";A 118");		//(assert (= (bv-or (bv-not (bv-redor (bool-to-bv (bv-gt #rx  #m )))) (bv-comp #B  0b1))   0b1)) ;118 BR
                                                    B <= #1 1'b1; $display(";A 120");		//(assert (= @B    0b1)) ;120 NB
                                                end
                                                else begin
                                                    $display(";A 119");		//(assert (= (bv-or (bv-not (bv-redor (bool-to-bv (bv-gt #rx  #m )))) (bv-comp #B  0b1))   0b0)) ;119 BR
                                                    B <= #1 1'b0; $display(";A 121");		//(assert (= @B    0b0)) ;121 NB
                                                end
                                            end
                                        4'b1101 :
                                            begin
                                                $display(";A 122");		//(assert (= #ff    0b1101)) ;122 CS
                                                if (((rx > m) || (B == 1'b1))) begin
                                                    $display(";A 123");		//(assert (= (bv-or (bool-to-bv (bv-gt #rx  #m )) (bv-comp #B  0b1))   0b1)) ;123 BR
                                                    B <= #1 1'b1; $display(";A 125");		//(assert (= @B    0b1)) ;125 NB
                                                end
                                                else begin
                                                    $display(";A 124");		//(assert (= (bv-or (bool-to-bv (bv-gt #rx  #m )) (bv-comp #B  0b1))   0b0)) ;124 BR
                                                    B <= #1 1'b0; $display(";A 126");		//(assert (= @B    0b0)) ;126 NB
                                                end
                                            end
                                        4'b1110 :
                                            begin
                                                $display(";A 127");		//(assert (= #ff    0b1110)) ;127 CS
                                                if ((rx > 31'b0111111111111111111111111111111)) begin
                                                    $display(";A 128");		//(assert (= (bool-to-bv (bv-gt #rx  0b0111111111111111111111111111111))   0b1)) ;128 BR
                                                    rx = rx; $display(";A 130");		//(assert (= @rx    #rx )) ;130 BL
                                                end
                                                else begin
                                                    $display(";A 129");		//(assert (= (bool-to-bv (bv-gt #rx  0b0111111111111111111111111111111))   0b0)) ;129 BR
                                                end
                                                if (((rx < m) || (B == 1'b1))) begin
                                                    $display(";A 131");		//(assert (= (bv-or (bool-to-bv (bv-lt #rx  #m )) (bv-comp #B  0b1))   0b1)) ;131 BR
                                                    B <= #1 1'b1; $display(";A 133");		//(assert (= @B    0b1)) ;133 NB
                                                end
                                                else begin
                                                    $display(";A 132");		//(assert (= (bv-or (bool-to-bv (bv-lt #rx  #m )) (bv-comp #B  0b1))   0b0)) ;132 BR
                                                    B <= #1 1'b0; $display(";A 134");		//(assert (= @B    0b0)) ;134 NB
                                                end
                                            end
                                        4'b1111 :
                                            begin
                                                $display(";A 135");		//(assert (= #ff    0b1111)) ;135 CS
                                                if ((rx > 31'b0111111111111111111111111111111)) begin
                                                    $display(";A 136");		//(assert (= (bool-to-bv (bv-gt #rx  0b0111111111111111111111111111111))   0b1)) ;136 BR
                                                    rx = rx; $display(";A 138");		//(assert (= @rx    #rx )) ;138 BL
                                                end
                                                else begin
                                                    $display(";A 137");		//(assert (= (bool-to-bv (bv-gt #rx  0b0111111111111111111111111111111))   0b0)) ;137 BR
                                                end
                                                if (((!(rx < m)) || (B == 1'b1))) begin
                                                    $display(";A 139");		//(assert (= (bv-or (bv-not (bv-redor (bool-to-bv (bv-lt #rx  #m )))) (bv-comp #B  0b1))   0b1)) ;139 BR
                                                    B <= #1 1'b1; $display(";A 141");		//(assert (= @B    0b1)) ;141 NB
                                                end
                                                else begin
                                                    $display(";A 140");		//(assert (= (bv-or (bv-not (bv-redor (bool-to-bv (bv-lt #rx  #m )))) (bv-comp #B  0b1))   0b0)) ;140 BR
                                                    B <= #1 1'b0; $display(";A 142");		//(assert (= @B    0b0)) ;142 NB
                                                end
                                            end
                                    endcase
                                end
                            1'b0 :
                                begin
                                    $display(";A 143");		//(assert (= #cf    0b0)) ;143 CS
                                    if ((df != 3'b111)) begin
                                        $display(";A 144");		//(assert (= (bv-not (bv-comp #df  0b111))   0b1)) ;144 BR
                                        if ((((df == 3'b101) && (B == 1'b0)) || ((df == 3'b100) && (B == 1'b1)))) begin
                                            $display(";A 146");		//(assert (= (bv-or (bv-and (bv-comp #df  0b101) (bv-comp #B  0b0)) (bv-and (bv-comp #df  0b100) (bv-comp #B  0b1)))   0b1)) ;146 BR
                                            d = 2'b11; $display(";A 148");		//(assert (= @d    0b11)) ;148 BL
                                        end
                                        else begin
                                            $display(";A 147");		//(assert (= (bv-or (bv-and (bv-comp #df  0b101) (bv-comp #B  0b0)) (bv-and (bv-comp #df  0b100) (bv-comp #B  0b1)))   0b0)) ;147 BR
                                            d = df[1:0]; $display(";A 149");		//(assert (= @d    (bv-extract 1 0 #df ))) ;149 BL
                                        end
                                        case (ff)
                                            4'b0000 :
                                                begin
                                                    $display(";A 150");		//(assert (= #ff    0b0000)) ;150 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 151");		//(assert (= #mf    0b00)) ;151 CS
                                                                m = {11'b00000000000, tail}; $display(";A 152");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;152 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 153");		//(assert (= #mf    0b01)) ;153 CS
                                                                m = datai; $display(";A 154");		//(assert (= @m    #datai )) ;154 BL
                                                                addr <= #1 tail; $display(";A 155");		//(assert (= @addr    #tail )) ;155 NB
                                                                rd <= #1 1'b1; $display(";A 156");		//(assert (= @rd    0b1)) ;156 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 157");		//(assert (= #mf    0b10)) ;157 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 158");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;158 NB
                                                                rd <= #1 1'b1; $display(";A 159");		//(assert (= @rd    0b1)) ;159 NB
                                                                m = datai; $display(";A 160");		//(assert (= @m    #datai )) ;160 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 161");		//(assert (= #mf    0b11)) ;161 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 162");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;162 NB
                                                                rd <= #1 1'b1; $display(";A 163");		//(assert (= @rd    0b1)) ;163 NB
                                                                m = datai; $display(";A 164");		//(assert (= @m    #datai )) ;164 BL
                                                            end
                                                    endcase
                                                    t = 31'b0000000000000000000000000000000; $display(";A 165");		//(assert (= @t    0b0000000000000000000000000000000)) ;165 BL
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 166");		//(assert (= #d    0b00)) ;166 CS
                                                                reg0 = (t - m); $display(";A 167");		//(assert (= @reg0    (bv-sub #t  #m ))) ;167 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 168");		//(assert (= #d    0b01)) ;168 CS
                                                                reg1 = (t - m); $display(";A 169");		//(assert (= @reg1    (bv-sub #t  #m ))) ;169 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 170");		//(assert (= #d    0b10)) ;170 CS
                                                                reg2 = (t - m); $display(";A 171");		//(assert (= @reg2    (bv-sub #t  #m ))) ;171 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 172");		//(assert (= #d    0b11)) ;172 CS
                                                                reg3 = (t - m); $display(";A 173");		//(assert (= @reg3    (bv-sub #t  #m ))) ;173 BL
                                                            end
                                                    endcase
                                                end
                                            4'b0001 :
                                                begin
                                                    $display(";A 174");		//(assert (= #ff    0b0001)) ;174 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 175");		//(assert (= #mf    0b00)) ;175 CS
                                                                m = {11'b00000000000, tail}; $display(";A 176");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;176 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 177");		//(assert (= #mf    0b01)) ;177 CS
                                                                m = datai; $display(";A 178");		//(assert (= @m    #datai )) ;178 BL
                                                                addr <= #1 tail; $display(";A 179");		//(assert (= @addr    #tail )) ;179 NB
                                                                rd <= #1 1'b1; $display(";A 180");		//(assert (= @rd    0b1)) ;180 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 181");		//(assert (= #mf    0b10)) ;181 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 182");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;182 NB
                                                                rd <= #1 1'b1; $display(";A 183");		//(assert (= @rd    0b1)) ;183 NB
                                                                m = datai; $display(";A 184");		//(assert (= @m    #datai )) ;184 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 185");		//(assert (= #mf    0b11)) ;185 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 186");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;186 NB
                                                                rd <= #1 1'b1; $display(";A 187");		//(assert (= @rd    0b1)) ;187 NB
                                                                m = datai; $display(";A 188");		//(assert (= @m    #datai )) ;188 BL
                                                            end
                                                    endcase
                                                    reg2 = reg3; $display(";A 189");		//(assert (= @reg2    #reg3 )) ;189 BL
                                                    reg3 = m; $display(";A 190");		//(assert (= @reg3    #m )) ;190 BL
                                                end
                                            4'b0010 :
                                                begin
                                                    $display(";A 191");		//(assert (= #ff    0b0010)) ;191 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 192");		//(assert (= #mf    0b00)) ;192 CS
                                                                m = {11'b00000000000, tail}; $display(";A 193");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;193 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 194");		//(assert (= #mf    0b01)) ;194 CS
                                                                m = datai; $display(";A 195");		//(assert (= @m    #datai )) ;195 BL
                                                                addr <= #1 tail; $display(";A 196");		//(assert (= @addr    #tail )) ;196 NB
                                                                rd <= #1 1'b1; $display(";A 197");		//(assert (= @rd    0b1)) ;197 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 198");		//(assert (= #mf    0b10)) ;198 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 199");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;199 NB
                                                                rd <= #1 1'b1; $display(";A 200");		//(assert (= @rd    0b1)) ;200 NB
                                                                m = datai; $display(";A 201");		//(assert (= @m    #datai )) ;201 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 202");		//(assert (= #mf    0b11)) ;202 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 203");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;203 NB
                                                                rd <= #1 1'b1; $display(";A 204");		//(assert (= @rd    0b1)) ;204 NB
                                                                m = datai; $display(";A 205");		//(assert (= @m    #datai )) ;205 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 206");		//(assert (= #d    0b00)) ;206 CS
                                                                reg0 = m; $display(";A 207");		//(assert (= @reg0    #m )) ;207 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 208");		//(assert (= #d    0b01)) ;208 CS
                                                                reg1 = m; $display(";A 209");		//(assert (= @reg1    #m )) ;209 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 210");		//(assert (= #d    0b10)) ;210 CS
                                                                reg2 = m; $display(";A 211");		//(assert (= @reg2    #m )) ;211 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 212");		//(assert (= #d    0b11)) ;212 CS
                                                                reg3 = m; $display(";A 213");		//(assert (= @reg3    #m )) ;213 BL
                                                            end
                                                    endcase
                                                end
                                            4'b0011 :
                                                begin
                                                    $display(";A 214");		//(assert (= #ff    0b0011)) ;214 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 215");		//(assert (= #mf    0b00)) ;215 CS
                                                                m = {11'b00000000000, tail}; $display(";A 216");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;216 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 217");		//(assert (= #mf    0b01)) ;217 CS
                                                                m = datai; $display(";A 218");		//(assert (= @m    #datai )) ;218 BL
                                                                addr <= #1 tail; $display(";A 219");		//(assert (= @addr    #tail )) ;219 NB
                                                                rd <= #1 1'b1; $display(";A 220");		//(assert (= @rd    0b1)) ;220 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 221");		//(assert (= #mf    0b10)) ;221 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 222");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;222 NB
                                                                rd <= #1 1'b1; $display(";A 223");		//(assert (= @rd    0b1)) ;223 NB
                                                                m = datai; $display(";A 224");		//(assert (= @m    #datai )) ;224 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 225");		//(assert (= #mf    0b11)) ;225 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 226");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;226 NB
                                                                rd <= #1 1'b1; $display(";A 227");		//(assert (= @rd    0b1)) ;227 NB
                                                                m = datai; $display(";A 228");		//(assert (= @m    #datai )) ;228 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 229");		//(assert (= #d    0b00)) ;229 CS
                                                                reg0 = m; $display(";A 230");		//(assert (= @reg0    #m )) ;230 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 231");		//(assert (= #d    0b01)) ;231 CS
                                                                reg1 = m; $display(";A 232");		//(assert (= @reg1    #m )) ;232 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 233");		//(assert (= #d    0b10)) ;233 CS
                                                                reg2 = m; $display(";A 234");		//(assert (= @reg2    #m )) ;234 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 235");		//(assert (= #d    0b11)) ;235 CS
                                                                reg3 = m; $display(";A 236");		//(assert (= @reg3    #m )) ;236 BL
                                                            end
                                                    endcase
                                                end
                                            4'b0100 :
                                                begin
                                                    $display(";A 237");		//(assert (= #ff    0b0100)) ;237 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 238");		//(assert (= #mf    0b00)) ;238 CS
                                                                m = {11'b00000000000, tail}; $display(";A 239");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;239 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 240");		//(assert (= #mf    0b01)) ;240 CS
                                                                m = datai; $display(";A 241");		//(assert (= @m    #datai )) ;241 BL
                                                                addr <= #1 tail; $display(";A 242");		//(assert (= @addr    #tail )) ;242 NB
                                                                rd <= #1 1'b1; $display(";A 243");		//(assert (= @rd    0b1)) ;243 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 244");		//(assert (= #mf    0b10)) ;244 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 245");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;245 NB
                                                                rd <= #1 1'b1; $display(";A 246");		//(assert (= @rd    0b1)) ;246 NB
                                                                m = datai; $display(";A 247");		//(assert (= @m    #datai )) ;247 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 248");		//(assert (= #mf    0b11)) ;248 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 249");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;249 NB
                                                                rd <= #1 1'b1; $display(";A 250");		//(assert (= @rd    0b1)) ;250 NB
                                                                m = datai; $display(";A 251");		//(assert (= @m    #datai )) ;251 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 252");		//(assert (= #d    0b00)) ;252 CS
                                                                reg0 = (rx + m); $display(";A 253");		//(assert (= @reg0    (bv-add #rx  #m ))) ;253 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 254");		//(assert (= #d    0b01)) ;254 CS
                                                                reg1 = (rx + m); $display(";A 255");		//(assert (= @reg1    (bv-add #rx  #m ))) ;255 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 256");		//(assert (= #d    0b10)) ;256 CS
                                                                reg2 = (rx + m); $display(";A 257");		//(assert (= @reg2    (bv-add #rx  #m ))) ;257 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 258");		//(assert (= #d    0b11)) ;258 CS
                                                                reg3 = (rx + m); $display(";A 259");		//(assert (= @reg3    (bv-add #rx  #m ))) ;259 BL
                                                            end
                                                    endcase
                                                end
                                            4'b0101 :
                                                begin
                                                    $display(";A 260");		//(assert (= #ff    0b0101)) ;260 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 261");		//(assert (= #mf    0b00)) ;261 CS
                                                                m = {11'b00000000000, tail}; $display(";A 262");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;262 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 263");		//(assert (= #mf    0b01)) ;263 CS
                                                                m = datai; $display(";A 264");		//(assert (= @m    #datai )) ;264 BL
                                                                addr <= #1 tail; $display(";A 265");		//(assert (= @addr    #tail )) ;265 NB
                                                                rd <= #1 1'b1; $display(";A 266");		//(assert (= @rd    0b1)) ;266 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 267");		//(assert (= #mf    0b10)) ;267 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 268");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;268 NB
                                                                rd <= #1 1'b1; $display(";A 269");		//(assert (= @rd    0b1)) ;269 NB
                                                                m = datai; $display(";A 270");		//(assert (= @m    #datai )) ;270 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 271");		//(assert (= #mf    0b11)) ;271 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 272");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;272 NB
                                                                rd <= #1 1'b1; $display(";A 273");		//(assert (= @rd    0b1)) ;273 NB
                                                                m = datai; $display(";A 274");		//(assert (= @m    #datai )) ;274 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 275");		//(assert (= #d    0b00)) ;275 CS
                                                                reg0 = (rx + m); $display(";A 276");		//(assert (= @reg0    (bv-add #rx  #m ))) ;276 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 277");		//(assert (= #d    0b01)) ;277 CS
                                                                reg1 = (rx + m); $display(";A 278");		//(assert (= @reg1    (bv-add #rx  #m ))) ;278 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 279");		//(assert (= #d    0b10)) ;279 CS
                                                                reg2 = (rx + m); $display(";A 280");		//(assert (= @reg2    (bv-add #rx  #m ))) ;280 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 281");		//(assert (= #d    0b11)) ;281 CS
                                                                reg3 = (rx + m); $display(";A 282");		//(assert (= @reg3    (bv-add #rx  #m ))) ;282 BL
                                                            end
                                                    endcase
                                                end
                                            4'b0110 :
                                                begin
                                                    $display(";A 283");		//(assert (= #ff    0b0110)) ;283 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 284");		//(assert (= #mf    0b00)) ;284 CS
                                                                m = {11'b00000000000, tail}; $display(";A 285");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;285 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 286");		//(assert (= #mf    0b01)) ;286 CS
                                                                m = datai; $display(";A 287");		//(assert (= @m    #datai )) ;287 BL
                                                                addr <= #1 tail; $display(";A 288");		//(assert (= @addr    #tail )) ;288 NB
                                                                rd <= #1 1'b1; $display(";A 289");		//(assert (= @rd    0b1)) ;289 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 290");		//(assert (= #mf    0b10)) ;290 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 291");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;291 NB
                                                                rd <= #1 1'b1; $display(";A 292");		//(assert (= @rd    0b1)) ;292 NB
                                                                m = datai; $display(";A 293");		//(assert (= @m    #datai )) ;293 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 294");		//(assert (= #mf    0b11)) ;294 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 295");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;295 NB
                                                                rd <= #1 1'b1; $display(";A 296");		//(assert (= @rd    0b1)) ;296 NB
                                                                m = datai; $display(";A 297");		//(assert (= @m    #datai )) ;297 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 298");		//(assert (= #d    0b00)) ;298 CS
                                                                reg0 = (rx - m); $display(";A 299");		//(assert (= @reg0    (bv-sub #rx  #m ))) ;299 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 300");		//(assert (= #d    0b01)) ;300 CS
                                                                reg1 = (rx - m); $display(";A 301");		//(assert (= @reg1    (bv-sub #rx  #m ))) ;301 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 302");		//(assert (= #d    0b10)) ;302 CS
                                                                reg2 = (rx - m); $display(";A 303");		//(assert (= @reg2    (bv-sub #rx  #m ))) ;303 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 304");		//(assert (= #d    0b11)) ;304 CS
                                                                reg3 = (rx - m); $display(";A 305");		//(assert (= @reg3    (bv-sub #rx  #m ))) ;305 BL
                                                            end
                                                    endcase
                                                end
                                            4'b0111 :
                                                begin
                                                    $display(";A 306");		//(assert (= #ff    0b0111)) ;306 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 307");		//(assert (= #mf    0b00)) ;307 CS
                                                                m = {11'b00000000000, tail}; $display(";A 308");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;308 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 309");		//(assert (= #mf    0b01)) ;309 CS
                                                                m = datai; $display(";A 310");		//(assert (= @m    #datai )) ;310 BL
                                                                addr <= #1 tail; $display(";A 311");		//(assert (= @addr    #tail )) ;311 NB
                                                                rd <= #1 1'b1; $display(";A 312");		//(assert (= @rd    0b1)) ;312 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 313");		//(assert (= #mf    0b10)) ;313 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 314");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;314 NB
                                                                rd <= #1 1'b1; $display(";A 315");		//(assert (= @rd    0b1)) ;315 NB
                                                                m = datai; $display(";A 316");		//(assert (= @m    #datai )) ;316 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 317");		//(assert (= #mf    0b11)) ;317 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 318");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;318 NB
                                                                rd <= #1 1'b1; $display(";A 319");		//(assert (= @rd    0b1)) ;319 NB
                                                                m = datai; $display(";A 320");		//(assert (= @m    #datai )) ;320 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 321");		//(assert (= #d    0b00)) ;321 CS
                                                                reg0 = (rx - m); $display(";A 322");		//(assert (= @reg0    (bv-sub #rx  #m ))) ;322 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 323");		//(assert (= #d    0b01)) ;323 CS
                                                                reg1 = (rx - m); $display(";A 324");		//(assert (= @reg1    (bv-sub #rx  #m ))) ;324 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 325");		//(assert (= #d    0b10)) ;325 CS
                                                                reg2 = (rx - m); $display(";A 326");		//(assert (= @reg2    (bv-sub #rx  #m ))) ;326 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 327");		//(assert (= #d    0b11)) ;327 CS
                                                                reg3 = (rx - m); $display(";A 328");		//(assert (= @reg3    (bv-sub #rx  #m ))) ;328 BL
                                                            end
                                                    endcase
                                                end
                                            4'b1000 :
                                                begin
                                                    $display(";A 329");		//(assert (= #ff    0b1000)) ;329 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 330");		//(assert (= #mf    0b00)) ;330 CS
                                                                m = {11'b00000000000, tail}; $display(";A 331");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;331 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 332");		//(assert (= #mf    0b01)) ;332 CS
                                                                m = datai; $display(";A 333");		//(assert (= @m    #datai )) ;333 BL
                                                                addr <= #1 tail; $display(";A 334");		//(assert (= @addr    #tail )) ;334 NB
                                                                rd <= #1 1'b1; $display(";A 335");		//(assert (= @rd    0b1)) ;335 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 336");		//(assert (= #mf    0b10)) ;336 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 337");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;337 NB
                                                                rd <= #1 1'b1; $display(";A 338");		//(assert (= @rd    0b1)) ;338 NB
                                                                m = datai; $display(";A 339");		//(assert (= @m    #datai )) ;339 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 340");		//(assert (= #mf    0b11)) ;340 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 341");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;341 NB
                                                                rd <= #1 1'b1; $display(";A 342");		//(assert (= @rd    0b1)) ;342 NB
                                                                m = datai; $display(";A 343");		//(assert (= @m    #datai )) ;343 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 344");		//(assert (= #d    0b00)) ;344 CS
                                                                reg0 = (rx + m); $display(";A 345");		//(assert (= @reg0    (bv-add #rx  #m ))) ;345 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 346");		//(assert (= #d    0b01)) ;346 CS
                                                                reg1 = (rx + m); $display(";A 347");		//(assert (= @reg1    (bv-add #rx  #m ))) ;347 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 348");		//(assert (= #d    0b10)) ;348 CS
                                                                reg2 = (rx + m); $display(";A 349");		//(assert (= @reg2    (bv-add #rx  #m ))) ;349 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 350");		//(assert (= #d    0b11)) ;350 CS
                                                                reg3 = (rx + m); $display(";A 351");		//(assert (= @reg3    (bv-add #rx  #m ))) ;351 BL
                                                            end
                                                    endcase
                                                end
                                            4'b1001 :
                                                begin
                                                    $display(";A 352");		//(assert (= #ff    0b1001)) ;352 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 353");		//(assert (= #mf    0b00)) ;353 CS
                                                                m = {11'b00000000000, tail}; $display(";A 354");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;354 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 355");		//(assert (= #mf    0b01)) ;355 CS
                                                                m = datai; $display(";A 356");		//(assert (= @m    #datai )) ;356 BL
                                                                addr <= #1 tail; $display(";A 357");		//(assert (= @addr    #tail )) ;357 NB
                                                                rd <= #1 1'b1; $display(";A 358");		//(assert (= @rd    0b1)) ;358 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 359");		//(assert (= #mf    0b10)) ;359 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 360");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;360 NB
                                                                rd <= #1 1'b1; $display(";A 361");		//(assert (= @rd    0b1)) ;361 NB
                                                                m = datai; $display(";A 362");		//(assert (= @m    #datai )) ;362 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 363");		//(assert (= #mf    0b11)) ;363 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 364");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;364 NB
                                                                rd <= #1 1'b1; $display(";A 365");		//(assert (= @rd    0b1)) ;365 NB
                                                                m = datai; $display(";A 366");		//(assert (= @m    #datai )) ;366 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 367");		//(assert (= #d    0b00)) ;367 CS
                                                                reg0 = (rx - m); $display(";A 368");		//(assert (= @reg0    (bv-sub #rx  #m ))) ;368 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 369");		//(assert (= #d    0b01)) ;369 CS
                                                                reg1 = (rx - m); $display(";A 370");		//(assert (= @reg1    (bv-sub #rx  #m ))) ;370 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 371");		//(assert (= #d    0b10)) ;371 CS
                                                                reg2 = (rx - m); $display(";A 372");		//(assert (= @reg2    (bv-sub #rx  #m ))) ;372 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 373");		//(assert (= #d    0b11)) ;373 CS
                                                                reg3 = (rx - m); $display(";A 374");		//(assert (= @reg3    (bv-sub #rx  #m ))) ;374 BL
                                                            end
                                                    endcase
                                                end
                                            4'b1010 :
                                                begin
                                                    $display(";A 375");		//(assert (= #ff    0b1010)) ;375 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 376");		//(assert (= #mf    0b00)) ;376 CS
                                                                m = {11'b00000000000, tail}; $display(";A 377");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;377 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 378");		//(assert (= #mf    0b01)) ;378 CS
                                                                m = datai; $display(";A 379");		//(assert (= @m    #datai )) ;379 BL
                                                                addr <= #1 tail; $display(";A 380");		//(assert (= @addr    #tail )) ;380 NB
                                                                rd <= #1 1'b1; $display(";A 381");		//(assert (= @rd    0b1)) ;381 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 382");		//(assert (= #mf    0b10)) ;382 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 383");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;383 NB
                                                                rd <= #1 1'b1; $display(";A 384");		//(assert (= @rd    0b1)) ;384 NB
                                                                m = datai; $display(";A 385");		//(assert (= @m    #datai )) ;385 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 386");		//(assert (= #mf    0b11)) ;386 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 387");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;387 NB
                                                                rd <= #1 1'b1; $display(";A 388");		//(assert (= @rd    0b1)) ;388 NB
                                                                m = datai; $display(";A 389");		//(assert (= @m    #datai )) ;389 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 390");		//(assert (= #d    0b00)) ;390 CS
                                                                reg0 = (rx + m); $display(";A 391");		//(assert (= @reg0    (bv-add #rx  #m ))) ;391 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 392");		//(assert (= #d    0b01)) ;392 CS
                                                                reg1 = (rx + m); $display(";A 393");		//(assert (= @reg1    (bv-add #rx  #m ))) ;393 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 394");		//(assert (= #d    0b10)) ;394 CS
                                                                reg2 = (rx + m); $display(";A 395");		//(assert (= @reg2    (bv-add #rx  #m ))) ;395 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 396");		//(assert (= #d    0b11)) ;396 CS
                                                                reg3 = (rx + m); $display(";A 397");		//(assert (= @reg3    (bv-add #rx  #m ))) ;397 BL
                                                            end
                                                    endcase
                                                end
                                            4'b1011 :
                                                begin
                                                    $display(";A 398");		//(assert (= #ff    0b1011)) ;398 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 399");		//(assert (= #mf    0b00)) ;399 CS
                                                                m = {11'b00000000000, tail}; $display(";A 400");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;400 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 401");		//(assert (= #mf    0b01)) ;401 CS
                                                                m = datai; $display(";A 402");		//(assert (= @m    #datai )) ;402 BL
                                                                addr <= #1 tail; $display(";A 403");		//(assert (= @addr    #tail )) ;403 NB
                                                                rd <= #1 1'b1; $display(";A 404");		//(assert (= @rd    0b1)) ;404 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 405");		//(assert (= #mf    0b10)) ;405 CS
                                                                addr <= #1 (tail + reg1[19:0]); $display(";A 406");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg1 )))) ;406 NB
                                                                rd <= #1 1'b1; $display(";A 407");		//(assert (= @rd    0b1)) ;407 NB
                                                                m = datai; $display(";A 408");		//(assert (= @m    #datai )) ;408 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 409");		//(assert (= #mf    0b11)) ;409 CS
                                                                addr <= #1 (tail + reg2[19:0]); $display(";A 410");		//(assert (= @addr    (bv-add #tail  (bv-extract 19 0 #reg2 )))) ;410 NB
                                                                rd <= #1 1'b1; $display(";A 411");		//(assert (= @rd    0b1)) ;411 NB
                                                                m = datai; $display(";A 412");		//(assert (= @m    #datai )) ;412 BL
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 413");		//(assert (= #d    0b00)) ;413 CS
                                                                reg0 = (rx - m); $display(";A 414");		//(assert (= @reg0    (bv-sub #rx  #m ))) ;414 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 415");		//(assert (= #d    0b01)) ;415 CS
                                                                reg1 = (rx - m); $display(";A 416");		//(assert (= @reg1    (bv-sub #rx  #m ))) ;416 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 417");		//(assert (= #d    0b10)) ;417 CS
                                                                reg2 = (rx - m); $display(";A 418");		//(assert (= @reg2    (bv-sub #rx  #m ))) ;418 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 419");		//(assert (= #d    0b11)) ;419 CS
                                                                reg3 = (rx - m); $display(";A 420");		//(assert (= @reg3    (bv-sub #rx  #m ))) ;420 BL
                                                            end
                                                    endcase
                                                end
                                            4'b1100 :
                                                begin
                                                    $display(";A 421");		//(assert (= #ff    0b1100)) ;421 CS
                                                    case (mf)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 422");		//(assert (= #mf    0b00)) ;422 CS
                                                                t = {1'b0, rx[30:1]}; $display(";A 423");		//(assert (= @t    (bv-concat 0b0 (bv-extract 30 1 #rx )))) ;423 BL
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 424");		//(assert (= #mf    0b01)) ;424 CS
                                                                t = {1'b0, ((B == 1'b1) ? 1'b0 : rx[30]), rx[29:1]}; $display(";A 425");		//(assert (= @t    (bv-concat 0b0 (ite (= (bv-comp #B  0b1) 0b1) 0b0 (bv-extract 30 30 #rx )) (bv-extract 29 1 #rx )))) ;425 BL
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 426");		//(assert (= #mf    0b10)) ;426 CS
                                                                t = {rx[29:0], 1'b0}; $display(";A 427");		//(assert (= @t    (bv-concat (bv-extract 29 0 #rx ) 0b0))) ;427 BL
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 428");		//(assert (= #mf    0b11)) ;428 CS
                                                                t = {rx[29:0], 1'b0}; $display(";A 429");		//(assert (= @t    (bv-concat (bv-extract 29 0 #rx ) 0b0))) ;429 BL
                                                                if ((t > 31'b0111111111111111111111111111111)) begin
                                                                    $display(";A 430");		//(assert (= (bool-to-bv (bv-gt #t  0b0111111111111111111111111111111))   0b1)) ;430 BR
                                                                    B <= #1 1'b1; $display(";A 432");		//(assert (= @B    0b1)) ;432 NB
                                                                end
                                                                else begin
                                                                    $display(";A 431");		//(assert (= (bool-to-bv (bv-gt #t  0b0111111111111111111111111111111))   0b0)) ;431 BR
                                                                    B <= #1 1'b0; $display(";A 433");		//(assert (= @B    0b0)) ;433 NB
                                                                end
                                                            end
                                                    endcase
                                                    case (d)
                                                        2'b00 :
                                                            begin
                                                                $display(";A 434");		//(assert (= #d    0b00)) ;434 CS
                                                                reg0 <= #1 t; $display(";A 435");		//(assert (= @reg0    #t )) ;435 NB
                                                            end
                                                        2'b01 :
                                                            begin
                                                                $display(";A 436");		//(assert (= #d    0b01)) ;436 CS
                                                                reg1 <= #1 t; $display(";A 437");		//(assert (= @reg1    #t )) ;437 NB
                                                            end
                                                        2'b10 :
                                                            begin
                                                                $display(";A 438");		//(assert (= #d    0b10)) ;438 CS
                                                                reg2 <= #1 t; $display(";A 439");		//(assert (= @reg2    #t )) ;439 NB
                                                            end
                                                        2'b11 :
                                                            begin
                                                                $display(";A 440");		//(assert (= #d    0b11)) ;440 CS
                                                                reg3 <= #1 t; $display(";A 441");		//(assert (= @reg3    #t )) ;441 NB
                                                            end
                                                    endcase
                                                end
                                        endcase
                                    end
                                    else begin
                                        $display(";A 145");		//(assert (= (bv-not (bv-comp #df  0b111))   0b0)) ;145 BR
                                        if ((df == 3'b111)) begin
                                            $display(";A 442");		//(assert (= (bv-comp #df  0b111)   0b1)) ;442 BR
                                            case (mf)
                                                2'b00 :
                                                    begin
                                                        $display(";A 444");		//(assert (= #mf    0b00)) ;444 CS
                                                        m = {11'b00000000000, tail}; $display(";A 445");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;445 BL
                                                    end
                                                2'b01 :
                                                    begin
                                                        $display(";A 446");		//(assert (= #mf    0b01)) ;446 CS
                                                        m = {11'b00000000000, tail}; $display(";A 447");		//(assert (= @m    (bv-concat 0b00000000000 #tail ))) ;447 BL
                                                    end
                                                2'b10 :
                                                    begin
                                                        $display(";A 448");		//(assert (= #mf    0b10)) ;448 CS
                                                        m = (reg1 + {11'b00000000000, tail}); $display(";A 449");		//(assert (= @m    (bv-add #reg1  (bv-concat 0b00000000000 #tail )))) ;449 BL
                                                    end
                                                2'b11 :
                                                    begin
                                                        $display(";A 450");		//(assert (= #mf    0b11)) ;450 CS
                                                        m = (reg2 + {11'b00000000000, tail}); $display(";A 451");		//(assert (= @m    (bv-add #reg2  (bv-concat 0b00000000000 #tail )))) ;451 BL
                                                    end
                                            endcase
                                            addr <= #1 m[19:0]; $display(";A 452");		//(assert (= @addr    (bv-extract 19 0 #m ))) ;452 NB
                                            wr <= #1 1'b1; $display(";A 453");		//(assert (= @wr    0b1)) ;453 NB
                                            datao <= #1 rx; $display(";A 454");		//(assert (= @datao    #rx )) ;454 NB
                                        end
                                        else begin
                                            $display(";A 443");		//(assert (= (bv-comp #df  0b111)   0b0)) ;443 BR
                                        end
                                    end
                                end
                        endcase
                        state <= #1 1'b0; $display(";A 455");		//(assert (= @state    0b0)) ;455 NB
                    end
            endcase
        end
    end

endmodule

